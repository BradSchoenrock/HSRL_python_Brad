netcdf out {
dimensions:
	altitude = 0 ;
	bin_range = 0 ;
	calibration = UNLIMITED ; 
	sondenamelength = 6 ;
	githash = 40 ;
	i2header = 1000 ;
	apheader = 1000 ;
	geoheader = 1000 ;
variables:
	int base_time ;
		base_time:string = "2006-10-23 18:19:59 UTC" ;
		base_time:long_name = "Base seconds since Unix Epoch" ;
		base_time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		base_time:dpl_py_binding = "dne" ;
	double sonde_times(calibration) ;
		sonde_times:long_name = "Time of Temperature Profiles" ;
		sonde_times:description = "New raob data" ;
		sonde_times:dpl_py_binding = "sounding.times" ;
        sonde_times:dpl_py_type = "python_datetime" ;
	double sonde_longitude(calibration) ;
		sonde_longitude:long_name = "Longitude of Temperature Profiles" ;
		sonde_longitude:units = "degree_E" ;
		sonde_longitude:description = "Sounding Longitude source" ;
		sonde_longitude:dpl_py_binding = "sounding.longitude" ;
	double sonde_latitude(calibration) ;
		sonde_latitude:long_name = "Latituide of Temperature Profiles" ;
		sonde_latitude:units = "degree_N" ;
		sonde_latitude:description = "Sounding Latitude source" ;
		sonde_latitude:dpl_py_binding = "sounding.latitude" ;
	double new_cal_times(calibration) ;
		new_cal_times:long_name = "Time of Calibration Change" ;
		new_cal_times:description = "New raob or system calibration data triggered recalibration" ;
		new_cal_times:dpl_py_binding = "chunk_start_time" ;
        new_cal_times:dpl_py_type = "python_datetime" ;
	float altitude(altitude) ;
		altitude:long_name = "Height above lidar" ;
		altitude:units = "meters" ;
		altitude:dpl_py_binding = "rs_mean.msl_altitudes" ;
	char calibration_version(calibration, githash) ;
		calibration_version:long_name = "Calibration Tables GIT Version" ;
		calibration_version:dpl_py_binding = "gitversion" ;
	byte new_cal_trigger(calibration) ;
		new_cal_trigger:long_name = "Trigger of Calibration Change" ;
		new_cal_trigger:description = "reason for recalibration" ;
		new_cal_trigger:bit_0 = "radiosonde profile" ;
		new_cal_trigger:bit_1 = "i2 scan" ;
		new_cal_trigger:bit_2 = "geometry" ;
		new_cal_trigger:dpl_py_binding = "dne" ;
	short new_cal_offset(calibration) ;
		new_cal_offset:long_name = "Record Dimension equivalent Offset" ;
		new_cal_offset:min_value = 0 ;
		new_cal_offset:dpl_py_binding = "dne" ;
	float top_alt_sounding(calibration) ;
		top_alt_sounding:long_name = "Sounding Maximum Altitude" ;
		top_alt_sounding:units = "meters" ;
		top_alt_sounding:dpl_py_binding = "sounding.top" ;
	float temperature_profile(calibration, altitude) ;
		temperature_profile:long_name = "Raob Temperature Profile" ;
		temperature_profile:description = "Temperature interpolated to requested altitude resolution" ;
		temperature_profile:units = "degrees Kelvin" ;
		temperature_profile:dpl_py_binding = "sounding.temps" ;
	float pressure_profile(calibration, altitude) ;
		pressure_profile:long_name = "Raob pressure Profile" ;
		pressure_profile:description = "Pressure interpolated to requested altitude resolution" ;
		pressure_profile:units = "hectopascals" ;
		pressure_profile:dpl_py_binding = "sounding.pressures" ;
	float dewpoint_profile(calibration, altitude) ;
		dewpoint_profile:long_name = "Raob Dewpoint Temperature Profile" ;
		dewpoint_profile:description = "Dewpoint interpolated to requested altitude resolution" ;
		dewpoint_profile:units = "degrees Kelvin" ;
		dewpoint_profile:missing_value = 9.96920996838687e+36 ;
		dewpoint_profile:dpl_py_binding = "sounding.dew_points" ;
	float windspeed_profile(calibration, altitude) ;
		windspeed_profile:long_name = "Raob Wind Speed Profile" ;
		windspeed_profile:description = "Speeds interpolated to requested altitude resolution" ;
		windspeed_profile:units = "m/s" ;
		windspeed_profile:missing_value = 9.96920996838687e+36 ;
		windspeed_profile:dpl_py_binding = "sounding.wind_spd" ;
	float winddir_profile(calibration, altitude) ;
		winddir_profile:long_name = "Raob Wind Direction Profile" ;
		winddir_profile:description = "Directions interpolated to requested altitude resolution" ;
		winddir_profile:units = "degrees" ;
		winddir_profile:missing_value = 9.96920996838687e+36 ;
		winddir_profile:dpl_py_binding = "sounding.wind_dir" ;
	char raob_station(calibration, sondenamelength) ;
		raob_station:long_name = "Radiosonde Station ID" ;
		raob_station:dpl_py_binding = "sounding.sounding_id" ;
	char i2_txt_header(calibration, i2header) ;
		i2_txt_header:long_name = "i2_scan_file_text_info" ;
		i2_txt_header:description = "Contains name of file used to compute calibration" ;
		i2_txt_header:dpl_py_binding = "dne" ;
	char geo_txt_header(calibration, geoheader) ;
		geo_txt_header:long_name = "geometric_correction_file_txt_header." ;
		geo_txt_header:dpl_py_binding = "dne" ;
	char ap_txt_header(calibration, apheader) ;
		ap_txt_header:long_name = "afterpulse_correction_file_txt_header." ;
		ap_txt_header:dpl_py_binding = "dne" ;
	double raob_time_offset(calibration) ;
		raob_time_offset:units = "seconds" ;
		raob_time_offset:long_name = "Radiosonde Launch time offset" ;
		raob_time_offset:description = "Time after base time in seconds" ;
		raob_time_offset:dpl_py_binding = "dne" ;
	short raob_time_vector(calibration) ;
		raob_time_vector:long_name = "Radiosonde Launch time vector" ;
		raob_time_vector:description = "Time in [year month day hour min sec ms us] format" ;
		raob_time_vector:dpl_py_binding = "dne" ;
	float Cmc(calibration, altitude) ;
		Cmc:long_name = "Molecular in Combined Calibration" ;
		Cmc:dpl_py_binding = "rs_Cxx.Cmc" ;
	float Cmm(calibration, altitude) ;
		Cmm:long_name = "Molecular in Molecular Calibration" ;
		Cmm:dpl_py_binding = "rs_Cxx.Cmm" ;
	float Cmm_i2a(calibration, altitude) ;
		Cmm_i2a:long_name = "Molecular i2a in Molecular i2a Calibration" ;
		Cmm_i2a:dpl_py_binding = "rs_Cxx.Cmm_i2a" ;
	float Cam(calibration) ;
		Cam:long_name = "Aerosol in Molecular Calibration" ;
		Cam:dpl_py_binding = "rs_Cxx.Cam" ;
	float Cam_i2a(calibration) ;
		Cam_i2a:long_name = "Aerosol in Molecular i2a Calibration" ;
		Cam_i2a:dpl_py_binding = "rs_Cxx.Cam_i2a" ;
	float beta_m(calibration, altitude) ;
		beta_m:long_name = "Raob molecular (Rayleigh) scattering cross section per unit volume" ;
		beta_m:units = "1/meter" ;
		beta_m:plot_scale = "logarithmic" ;
		beta_m:dpl_py_binding = "rs_Cxx.beta_r" ;
	float combined_gain(calibration) ;
		combined_gain:long_name = "Combined Gain Factor" ;
		combined_gain:description = "Low Gain level * Factor ~ High Gain level" ;
		combined_gain:dpl_py_binding = "rs_constants.hi_to_low_combined_channel_gain_ratio" ;
	float combined_merge_threshhold(calibration) ;
		combined_merge_threshhold:long_name = "Combined Merge Threshhold" ;
		combined_merge_threshhold:dpl_py_binding = "rs_constants.combined_channel_merge_threshhold" ;
	float polarization_cross_talk(calibration) ;
		polarization_cross_talk:long_name = "Polarization Cross Talk" ;
		polarization_cross_talk:dpl_py_binding = "rs_constants.polarization_cross_talk" ;
	float wfov_to_combined_gain_ratio(calibration) ;
		wfov_to_combined_gain_ratio:long_name = "WFOV to Combined Gain" ;
		wfov_to_combined_gain_ratio:dpl_py_binding = "rs_constants.wfov_to_combined_gain_ratio" ;
	float combined_to_cross_pol_gain_ratio(calibration) ;
		combined_to_cross_pol_gain_ratio:long_name = "Combined to Cross Pol Gain" ;
		combined_to_cross_pol_gain_ratio:dpl_py_binding = "rs_constants.combined_to_cross_pol_gain_ratio" ;
	float molecular_to_wfov_gain_ratio(calibration) ;
		molecular_to_wfov_gain_ratio:long_name = "Molecular to WFOV Gain" ;
		molecular_to_wfov_gain_ratio:dpl_py_binding = "rs_constants.molecular_to_wfov_gain_ratio" ;
	float geo_cor(calibration, bin_range) ;
		geo_cor:long_name = "Overlap correction" ;
		geo_cor:description = "Geometric overlap correction in raw range bins" ;
		geo_cor:units = " " ;
		geo_cor:missing_value = 9.96920996838687e+36 ;
		geo_cor:plot_scale = "logarithmic" ;
		geo_cor:dpl_py_binding = "geo_corr" ;

// global attributes:
        :dpl_py_template = "hsrl_calibration.cdl" ;
        :dpl_py_template_version = 20140625 ;
		:time_zone = "UTC" ;
}
