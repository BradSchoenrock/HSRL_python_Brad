netcdf out {
dimensions:
	time = UNLIMITED ;
	altitude = 0 ;
	stationid = 15 ;
	soundingid = 15 ;
	soundingtype = 15 ;
variables:
	int base_time ;
		base_time:string = "2006-10-23 18:19:59 UTC" ;
		base_time:long_name = "Base seconds since Unix Epoch" ;
		base_time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		base_time:dpl_py_binding = "dne" ;
	double time(time) ;
		time:long_name = "Time" ;
		time:units = "seconds since 2006-10-23 18:19:59 UTC" ;
		time:dpl_py_binding = "times" ;
        time:dpl_py_type = "python_datetime" ;
	double expire_time(time) ;
		expire_time:long_name = "Time" ;
		expire_time:units = "seconds since 2006-10-23 18:19:59 UTC" ;
		expire_time:dpl_py_binding = "expire_time" ;
        expire_time:dpl_py_type = "python_datetime" ;
	float latitude(time) ;
		latitude:long_name = "latitude of lidar" ;
		latitude:units = "degree_N" ;
		latitude:dpl_py_binding = "latitude" ;
	float longitude(time) ;
		longitude:long_name = "longitude of lidar" ;
		longitude:units = "degree_E" ;
		longitude:dpl_py_binding = "longitude" ;
	float altitude(time,altitude) ;
		altitude:long_name = "Height above lidar" ;
		altitude:units = "meters" ;
		altitude:dpl_py_binding = "altitudes" ;
	float top_alt_sounding(time) ;
		top_alt_sounding:long_name = "Sounding Maximum Altitude" ;
		top_alt_sounding:units = "meters" ;
		top_alt_sounding:dpl_py_binding = "top" ;
	float bot_alt_sounding(time) ;
		bot_alt_sounding:long_name = "Sounding Minimum Altitude" ;
		bot_alt_sounding:units = "meters" ;
		bot_alt_sounding:dpl_py_binding = "bot" ;
	float temperature_profile(time, altitude) ;
		temperature_profile:long_name = "Temperature Profile" ;
		temperature_profile:description = "Temperature" ;
		temperature_profile:units = "degrees Kelvin" ;
		temperature_profile:dpl_py_binding = "temps" ;
	float pressure_profile(time, altitude) ;
		pressure_profile:long_name = "Pressure Profile" ;
		pressure_profile:description = "Pressure" ;
		pressure_profile:units = "hectopascals" ;
		pressure_profile:dpl_py_binding = "pressures" ;
	float dewpoint_profile(time, altitude) ;
		dewpoint_profile:long_name = "Dewpoint Temperature Profile" ;
		dewpoint_profile:description = "Dewpoint" ;
		dewpoint_profile:units = "degrees Kelvin" ;
		dewpoint_profile:missing_value = 9.96920996838687e+36 ;
		dewpoint_profile:dpl_py_binding = "dew_points" ;
	float frostpoint_profile(time, altitude) ;
		frostpoint_profile:long_name = "Frostpoint Temperature Profile" ;
		frostpoint_profile:description = "Frostpoint" ;
		frostpoint_profile:units = "degrees Kelvin" ;
		frostpoint_profile:missing_value = 9.96920996838687e+36 ;
		frostpoint_profile:dpl_py_binding = "frost_points" ;
	char station(time, stationid) ;
		station:long_name = "Radiosonde Station ID" ;
		station:dpl_py_binding = "station_id" ;
	char sounding(time, soundingid) ;
		sounding:long_name = "Radiosonde Station ID" ;
		sounding:dpl_py_binding = "sounding_id" ;
	char sounding_type(time,soundingtype) ;
		sounding_type:long_name = "Radiosonde Station ID" ;
		sounding_type:dpl_py_binding = "sounding_type" ;

// global attributes:
        :dpl_py_template = "NWS_Profile_Archive.cdl" ;
        :dpl_py_template_version = 20141001 ;
		:time_zone = "UTC" ;
}
