netcdf out {
dimensions:
	time = UNLIMITED ;
	altitude = 0 ;
	time_vector = 8 ;
variables:
	int base_time ;
		base_time:string = "2006-10-23 18:19:59 UTC" ;
		base_time:long_name = "Base seconds since Unix Epoch" ;
		base_time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		base_time:dpl_py_binding = "dne" ;
	short first_time(time_vector) ;
		first_time:long_name = "First Time in file" ;
		first_time:dpl_py_binding = "dne" ;
	short last_time(time_vector) ;
		last_time:long_name = "Last Time in file" ;
		last_time:dpl_py_binding = "dne" ;
	double time(time) ;
		time:long_name = "Time" ;
		time:units = "seconds since 2006-10-23 18:19:59 UTC" ;
		time:dpl_py_binding = "rs_inv.times" ;
                time:dpl_py_type = "python_datetime" ;
	double mean_time(time) ;
		mean_time:long_name = "Mean Time" ;
		mean_time:units = "seconds since 2006-10-23 18:19:59 UTC" ;
		mean_time:dpl_py_binding = "rs_mean.times" ;
        mean_time:dpl_py_type = "python_datetime" ;
	double time_offset(time) ;
		time_offset:long_name = "Time offset from base_time" ;
		time_offset:description = "same times as \"First time in record\" " ;
		time_offset:units = "seconds since 2006-10-23 18:19:59 UTC" ;
		time_offset:dpl_py_binding = "dne" ;
	short start_time(time, time_vector) ;
		start_time:long_name = "First Time in record" ;
		start_time:description = "time of first laser shot in averaging interval" ;
		start_time:dpl_py_binding = "dne" ;
	float latitude(time) ;
		latitude:long_name = "latitude of lidar" ;
		latitude:units = "degree_N" ;
		latitude:dpl_py_binding = "rs_mean.latitude" ;
	float longitude(time) ;
		longitude:long_name = "longitude of lidar" ;
		longitude:units = "degree_E" ;
		longitude:dpl_py_binding = "rs_mean.longitude" ;
	float lidar_altitude(time) ;
		lidar_altitude:long_name = "ground based platform altitude" ;
		lidar_altitude:units = "meters" ;
		lidar_altitude:dpl_py_binding = "rs_mean.GPS_MSL_Alt" ;
	float range_resolution ;
		range_resolution:long_name = "Range resolution" ;
		range_resolution:description = "vertical distance between data points after averaging" ;
		range_resolution:units = "meters" ;
		range_resolution:dpl_py_binding = "dne" ;
	float time_average ;
		time_average:long_name = "Time Averaging Width" ;
		time_average:description = "Time between data points after averaging" ;
		time_average:units = "seconds" ;
		time_average:dpl_py_binding = "dne" ;
	float transmitted_energy(time) ;
		transmitted_energy:long_name = "Transmitted Energy" ;
		transmitted_energy:units = "Joules" ;
		transmitted_energy:missing_value = 9.96920996838687e+36 ;
		transmitted_energy:dpl_py_binding = "rs_mean.transmitted_energy" ;
	float piezovoltage(time) ;
		piezovoltage:long_name = "piezovoltage" ;
		piezovoltage:units = "Volts" ;
		piezovoltage:missing_value = 9.96920996838687e+36 ;
		piezovoltage:dpl_py_binding = "dne" ;
	int num_seeded_shots(time) ;
		num_seeded_shots:long_name = "Number of Seeded Shots" ;
		num_seeded_shots:missing_value = -1 ;
		num_seeded_shots:dpl_py_binding = "rs_mean.seeded_shots" ;
	int num_shots(time) ;
		num_shots:long_name = "Number of Shots" ;
		num_shots:missing_value = -1 ;
		num_shots:dpl_py_binding = "rs_mean.shot_count" ;
	float seed_quality(time) ;
		seed_quality:long_name = "Laser Seeding Quality" ;
		seed_quality:description = "The ratio of seeded shots to total shots. Only seeded shot data is stored and processed.  A low seed ratio can result in low noise resistance." ;
		seed_quality:missing_value = 9.96920996838687e+36 ;
		seed_quality:range = 0., 1. ;
		seed_quality:dpl_py_binding = "dne" ;
	float frequency_quality(time) ;
		frequency_quality:long_name = "Laser Frequency Quality" ;
		frequency_quality:description = "An ratio average of how good the frequency lock is per raw interval. A low value can result in poor separation of molecular and aerosol counts." ;
		frequency_quality:missing_value = 9.96920996838687e+36 ;
		frequency_quality:range = 0., 1. ;
		frequency_quality:dpl_py_binding = "dne" ;
	float lock_quality(time) ;
		lock_quality:long_name = "Laser Lock Quality" ;
		lock_quality:description = "A ratio of likely locked intervals (frequency_quality>=.5) to seeded intervals.  A low value can result in poor separation of molecular and aerosol counts." ;
		lock_quality:missing_value = 9.96920996838687e+36 ;
		lock_quality:range = 0., 1. ;
		lock_quality:dpl_py_binding = "dne" ;
	float mol_cal_pulse(time) ;
		mol_cal_pulse:long_name = "Molecular calibration pulse" ;
		mol_cal_pulse:description = "Sum of photon counts in the molecular channel due to light scattered with the telescope." ;
		mol_cal_pulse:units = "counts" ;
		mol_cal_pulse:missing_value = 9.96920996838687e+36 ;
		mol_cal_pulse:dpl_py_binding = "rs_mean.molecular_cal_pulse" ;
	float mol_i2a_cal_pulse(time) ;
		mol_i2a_cal_pulse:long_name = "Molecular I2A calibration pulse" ;
		mol_i2a_cal_pulse:description = "Sum of photon counts in the molecular channel due to light scattered with the telescope." ;
		mol_i2a_cal_pulse:units = "counts" ;
		mol_i2a_cal_pulse:missing_value = 9.96920996838687e+36 ;
		mol_i2a_cal_pulse:dpl_py_binding = "rs_mean.molecular_i2a_cal_pulse" ;
	int mol_norm_idx ;
		mol_norm_idx:dpl_py_binding = "rs_inv.mol_norm_index" ;
	float c_pol_dark_count(time) ;
		c_pol_dark_count:long_name = "Cross Polarization Dark Count FIXME dark counts need alt" ;
		c_pol_dark_count:description = "total counts per averaging interval(eg. one altitude, one time)" ;
		c_pol_dark_count:units = "counts" ;
		c_pol_dark_count:missing_value = 9.96920996838687e+36 ;
		c_pol_dark_count:dpl_py_binding = "rs_mean.c_pol_dark_counts" ;
	float mol_i2a_dark_count(time) ;
		mol_i2a_dark_count:long_name = "Molecular I2A Dark Count" ;
		mol_i2a_dark_count:description = "total counts per averaging interval(eg. one altitude, one time)" ;
		mol_i2a_dark_count:units = "counts" ;
		mol_i2a_dark_count:missing_value = 9.96920996838687e+36 ;
		mol_i2a_dark_count:dpl_py_binding = "rs_mean.mol_i2a_dark_counts" ;
	float mol_dark_count(time) ;
		mol_dark_count:long_name = "Molecular Dark Count" ;
		mol_dark_count:description = "total counts per averaging interval(eg. one altitude, one time)" ;
		mol_dark_count:units = "counts" ;
		mol_dark_count:missing_value = 9.96920996838687e+36 ;
		mol_dark_count:dpl_py_binding = "rs_mean.mol_dark_counts" ;
	float combined_dark_count_lo(time) ;
		combined_dark_count_lo:long_name = "Low Gain Combined Dark Count" ;
		combined_dark_count_lo:description = "total counts per averaging interval(eg. one altitude, one time)" ;
		combined_dark_count_lo:units = "counts" ;
		combined_dark_count_lo:missing_value = 9.96920996838687e+36 ;
		combined_dark_count_lo:dpl_py_binding = "rs_mean.c_lo_dark_counts" ;
	float combined_dark_count_hi(time) ;
		combined_dark_count_hi:long_name = "High Gain Combined Dark Count" ;
		combined_dark_count_hi:description = "total counts per averaging interval(eg. one altitude, one time)" ;
		combined_dark_count_hi:units = "counts" ;
		combined_dark_count_hi:missing_value = 9.96920996838687e+36 ;
		combined_dark_count_hi:dpl_py_binding = "rs_mean.c_hi_dark_counts" ;
	int od_norm_index ;
		od_norm_index:long_name = "Optical depth normalization index FIXME shouldn't be needed" ;
		od_norm_index:dpl_py_binding = "rs_inv.od_norm_index" ;
	float od(time, altitude) ;
		od:long_name = "Optical depth of particulate" ;
		od:units = " " ;
		od:missing_value = 9.96920996838687e+36 ;
		od:insufficient_data = 9.96920996838687e+36 ;
		od:plot_scale = "logarithmic" ;
		od:dpl_py_binding = "rs_inv.optical_depth" ;
	float extinction(time,altitude) ;
		extinction:long_name = "Extinction Profile" ;
		extinction:units = " " ;
		extinction:missing_value = 9.96920996838687e+36 ;
		extinction:insufficient_data = 9.96920996838687e+36 ;
		extinction:plot_scale = "logarithmic" ;
		extinction:dpl_py_binding = "rs_inv.extinction" ;
	float effective_diameter_prime(time, altitude) ;
		effective_diameter_prime:long_name = "lidar/radar effective particle diameter" ;
		effective_diameter_prime:units = "microns" ;
		effective_diameter_prime:description = "Effective diameter directly from the ratio of Lidar Backscatter and Radar Reflectivity; (<volume^2>/<area>)^.25, see Donovan JGR Nov 2001" ;
		effective_diameter_prime:missing_value = 9.96920996838687e+36 ;
		effective_diameter_prime:dpl_py_binding = "dne" ;
	float effective_diameter(time, altitude) ;
		effective_diameter:long_name = "Effective particle diameter" ;
		effective_diameter:units = "microns" ;
		effective_diameter:description = "Effective particle diameter derived from ratio of Lidar Backscatter and Radar Reflectivity; assuming a gamma size distribution" ;
		effective_diameter:missing_value = 9.96920996838687e+36 ;
		effective_diameter:dpl_py_binding = "dne" ;
	float num_particles(time, altitude) ;
		num_particles:long_name = "Number density of particles" ;
		num_particles:units = "1/liter" ;
		num_particles:description = "Number of particles per liter derived from ratio of lidar backscatter and radar reflectivity; assuming a gamma size distribution" ;
		num_particles:missing_value = 9.96920996838687e+36 ;
		num_particles:dpl_py_binding = "dne" ;
	float mean_diameter(time, altitude) ;
		mean_diameter:long_name = "Mean diameter of particles" ;
		mean_diameter:units = "microns" ;
		mean_diameter:description = "Mean diameter of particles derived from the effective diameter and the gamma size distribution" ;
		mean_diameter:missing_value = 9.96920996838687e+36 ;
		mean_diameter:dpl_py_binding = "dne" ;
	float LWC(time, altitude) ;
		LWC:long_name = "Liquid water content" ;
		LWC:units = "gr/m^3" ;
		LWC:description = "Liquid water content derived from ratio of lidar backscatter and radar reflectivity; assuming a gamma size distribution" ;
		LWC:missing_value = 9.96920996838687e+36 ;
		LWC:dpl_py_binding = "dne" ;
	float beta_a(time, altitude) ;
		beta_a:long_name = "Particulate extinction cross section per unit volume" ;
		beta_a:units = "1/m" ;
		beta_a:missing_value = 9.96920996838687e+36 ;
		beta_a:plot_scale = "logarithmic" ;
		beta_a:dpl_py_binding = "dne" ;
	float atten_beta_r_backscat(time, altitude) ;
		atten_beta_r_backscat:long_name = "Attenuated Molecular return" ;
		atten_beta_r_backscat:units = "1/(m sr)" ;
		atten_beta_r_backscat:missing_value = 9.96920996838687e+36 ;
		atten_beta_r_backscat:plot_scale = "logarithmic" ;
		atten_beta_r_backscat:dpl_py_binding = "rs_inv.atten_beta_a_backscat" ;
	float circular_depol(time, altitude) ;
		circular_depol:long_name = "Circular depolarization ratio for particulate" ;
		circular_depol:description = "left circular return divided by right circular return" ;
		circular_depol:units = " " ;
		circular_depol:missing_value = 9.96920996838687e+36 ;
		circular_depol:plot_scale = "logarithmic" ;
		circular_depol:dpl_py_binding = "rs_inv.circular_depol" ;
	float linear_depol(time, altitude) ;
		linear_depol:long_name = "Linear depolarization ratio for particulate" ;
		linear_depol:description = "Linear depolarization return" ;
		linear_depol:units = " " ;
		linear_depol:missing_value = 9.96920996838687e+36 ;
		linear_depol:plot_scale = "logarithmic" ;
		linear_depol:dpl_py_binding = "rs_inv.linear_depol" ;
	float beta_a_backscat_parallel(time, altitude) ;
		beta_a_backscat_parallel:long_name = "Particulate nondepolarized backscatter cross section per unit volume" ;
		beta_a_backscat_parallel:units = "1/(m sr)" ;
		beta_a_backscat_parallel:missing_value = 9.96920996838687e+36 ;
		beta_a_backscat_parallel:plot_scale = "logarithmic" ;
		beta_a_backscat_parallel:dpl_py_binding = "rs_inv.beta_a_backscat_par" ;
	float beta_a_backscat(time, altitude) ;
		beta_a_backscat:long_name = "Particulate backscatter cross section per unit volume" ;
		beta_a_backscat:units = "1/(m sr)" ;
		beta_a_backscat:missing_value = 9.96920996838687e+36 ;
		beta_a_backscat:plot_scale = "logarithmic" ;
		beta_a_backscat:dpl_py_binding = "rs_inv.beta_a_backscat" ;
	float Na(time, altitude) ;
		Na:long_name = "Inverted Aerosol" ;
		Na:units = " " ;
		Na:dpl_py_binding = "rs_inv.Na" ;
	float Nm(time, altitude) ;
		Nm:long_name = "Inverted Molecular" ;
		Nm:units = " " ;
		Nm:dpl_py_binding = "rs_inv.Nm" ;
	float Nm_i2a(time, altitude) ;
		Nm_i2a:long_name = "Inverted I2A Molecular" ;
		Nm_i2a:units = " " ;
		Nm_i2a:dpl_py_binding = "rs_inv.Nm_i2a" ;
	float Ncp(time, altitude) ;
		Ncp:long_name = "Inverted Cross Polarization" ;
		Ncp:units = " " ;
		Ncp:dpl_py_binding = "rs_inv.Ncp" ;
	int qc_mask(time, altitude) ;
		qc_mask:long_name = "Quality Mask" ;
		qc_mask:description = "Quality mask bitfield.  Unused bits are always high" ;
		qc_mask:missing_value = 0 ;
		qc_mask:_Unsigned = "true" ;
		qc_mask:bit_0 = "complete_mask" ;
		qc_mask:bit_0_description = "data is good.  and of bits 1-9" ;
		qc_mask:bit_1 = "lidar_ok_mask" ;
		qc_mask:bit_1_description = "lidar data is present" ;
		qc_mask:bit_2 = "lock_quality_mask" ;
		qc_mask:bit_2_description = "laser is locked to iodine filter wavelength" ;
		qc_mask:bit_3 = "seed_quality_mask" ;
		qc_mask:bit_3_description = "laser wavelength is locked to seed laser" ;
		qc_mask:bit_4 = "mol_count_snr_mask" ;
		qc_mask:bit_4_description = "molecular signal/photon counting error in molecular signal is above specified threshhold" ;
		qc_mask:bit_5 = "backscat_snr_mask" ;
		qc_mask:bit_5_description = "backscatter cross-section/photon counting error in backscatter cross-section is above specified threshhold" ;
		qc_mask:bit_6 = "mol_lost_mask" ;
		qc_mask:bit_6_description = "number of molecular photon counts is above specified threshhold" ;
		qc_mask:bit_7 = "min_backscat_mask" ;
		qc_mask:bit_7_description = "lidar backscatter cross-section is above specified threshhold" ;
		qc_mask:bit_8 = "radar_backscat_mask" ;
		qc_mask:bit_8_description = "radar backscatter cross-section is above specified threshhold" ;
		qc_mask:bit_9 = "radar_ok_mask" ;
		qc_mask:bit_9_description = "radar data is present" ;
		qc_mask:bit_10 = "aeri_ok_mask" ;
		qc_mask:bit_10_description = "aeri data is present" ;
		qc_mask:bit_11 = "aeri_qc_mask" ;
		qc_mask:bit_11_description = "aeri data has passed a quality check" ;
		qc_mask:dpl_py_binding = "rs_inv.qc_mask" ;
	float std_beta_a_backscat(time, altitude) ;
		std_beta_a_backscat:long_name = "Std dev of backscat cross section (photon counting)" ;
		std_beta_a_backscat:units = "1/(m sr)" ;
		std_beta_a_backscat:missing_value = 9.96920996838687e+36 ;
		std_beta_a_backscat:plot_scale = "logarithmic" ;
		std_beta_a_backscat:dpl_py_binding = "dne" ;
	float mwr_frequency(mwr_frequency) ;
		mwr_frequency:long_name = "Frequency" ;
		mwr_frequency:units = "GHz" ;
		mwr_frequency:missing_value = 9.96920996838687e+36 ;
		mwr_frequency:dpl_py_binding = "dne" ;
	float mwr_btemp(time, mwr_frequency) ;
		mwr_btemp:long_name = "MWR Brightness Temperature" ;
		mwr_btemp:units = "degK" ;
		mwr_btemp:missing_value = 9.96920996838687e+36 ;
		mwr_btemp:dpl_py_binding = "dne" ;

// global attributes:
                :dpl_py_template = "segment_hsrl_processed.cdl" ;
                :dpl_py_template_version = 20140216 ;
		:time_zone = "UTC" ;
}
