netcdf out {
dimensions:
    time = UNLIMITED ;
    raw_time = UNLIMITED ;
    altitude = 0 ;
    bin_range = 0;
    profile_time = 1;
    time_vector = 8 ;
    calibration = UNLIMITED ; 
    sondenamelength = 32 ;
    githash = 40 ;
    i2header = 2000 ;
    geoheader = 2000 ;
    apheader = 2000 ;
    aeri_btemp_wavenumber = 0 ;
    aeri_mean_rad_wavenumber_ch1 = 0 ;
    aeri_mean_rad_wavenumber_ch2 = 0 ;
    mwr_frequency = 0 ;
    uncertainty = 2 ;
variables:
    int base_time ;
        base_time:string = "2006-10-23 18:19:59 UTC" ;
        base_time:long_name = "Base seconds since Unix Epoch" ;
        base_time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
        base_time:dpl_py_binding = "dne" ;
    short first_time(time_vector) ;
        first_time:long_name = "First Time in file" ;
        first_time:dpl_py_binding = "dne" ;
    short last_time(time_vector) ;
        last_time:long_name = "Last Time in file" ;
        last_time:dpl_py_binding = "dne" ;
    double time(time) ;
        time:long_name = "Time" ;
        time:units = "seconds since 2006-10-23 18:19:59 UTC" ;
        time:dpl_py_binding = "rs_inv.times" ;
        time:dpl_py_type = "python_datetime" ;
    double mean_time(time) ;
        mean_time:long_name = "Mean Time" ;
        mean_time:units = "seconds since 2006-10-23 18:19:59 UTC" ;
        mean_time:dpl_py_binding = "rs_mean.times" ;
        mean_time:dpl_py_type = "python_datetime" ;
    double raw_time(raw_time) ;
        raw_time:long_name = "Raw Time" ;
        raw_time:units = "seconds since 2006-10-23 18:19:59 UTC" ;
        raw_time:dpl_py_binding = "rs_raw.times" ;
        raw_time:dpl_py_type = "python_datetime" ;
    double time_offset(time) ;
        time_offset:long_name = "Time offset from base_time" ;
        time_offset:description = "same times as \"First time in record\" " ;
        time_offset:units = "seconds since 2006-10-23 18:19:59 UTC" ;
        time_offset:dpl_py_binding = "dne" ;
    short start_time(time, time_vector) ;
        start_time:long_name = "First Time in record" ;
        start_time:description = "time of first laser shot in averaging interval" ;
        start_time:dpl_py_binding = "dne" ;
    float latitude(time) ;
        latitude:long_name = "latitude of lidar" ;
        latitude:units = "degree_N" ;
        latitude:dpl_py_binding = "rs_mean.latitude" ;
    float longitude(time) ;
        longitude:long_name = "longitude of lidar" ;
        longitude:units = "degree_E" ;
        longitude:dpl_py_binding = "rs_mean.longitude" ;
    float telescope_roll_angle_offset(time) ;
        telescope_roll_angle_offset:long_name = "Telescope Mounting Roll Angle Offset" ;
        telescope_roll_angle_offset:description = "Telescope Mount Roll Angle Relative to aircraft up measured clockwise" ;
        telescope_roll_angle_offset:units = "degrees" ;
        telescope_roll_angle_offset:range = -180.0, 360.0 ;
        telescope_roll_angle_offset:dpl_py_binding = "rs_mean.telescope_roll_angle_offset" ;
    float lidar_altitude(time) ;
        lidar_altitude:long_name = "ground based platform altitude" ;
        lidar_altitude:units = "meters" ;
        lidar_altitude:dpl_py_binding = "rs_mean.GPS_MSL_Alt" ;
    float range_resolution ;
        range_resolution:long_name = "Range resolution" ;
        range_resolution:description = "vertical distance between data points after averaging" ;
        range_resolution:units = "meters" ;
        range_resolution:dpl_py_binding = "dne" ;
    float time_average ;
        time_average:long_name = "Time Averaging Width" ;
        time_average:description = "Time between data points after averaging" ;
        time_average:units = "seconds" ;
        time_average:dpl_py_binding = "dne" ;
    double sonde_times(calibration) ;
        sonde_times:long_name = "Time of Temperature Profiles" ;
        sonde_times:description = "New raob data" ;
        sonde_times:dpl_py_binding = "sounding.times" ;
        sonde_times:dpl_py_type = "python_datetime" ;
    double sonde_longitude(calibration) ;
        sonde_longitude:long_name = "Longitude of Temperature Profiles" ;
        sonde_longitude:units = "degree_E" ;
        sonde_longitude:description = "Sounding Longitude source" ;
        sonde_longitude:dpl_py_binding = "sounding.longitude" ;
    double sonde_latitude(calibration) ;
        sonde_latitude:long_name = "Latituide of Temperature Profiles" ;
        sonde_latitude:units = "degree_N" ;
        sonde_latitude:description = "Sounding Latitude source" ;
        sonde_latitude:dpl_py_binding = "sounding.latitude" ;
    double new_cal_times(calibration) ;
        new_cal_times:long_name = "Time of Calibration Change" ;
        new_cal_times:description = "New raob or system calibration data triggered recalibration" ;
        new_cal_times:dpl_py_binding = "chunk_start_time" ;
        new_cal_times:dpl_py_type = "python_datetime" ;
    float altitude(altitude) ;
        altitude:long_name = "Height above lidar" ;
        altitude:units = "meters" ;
        altitude:dpl_py_binding = "rs_mean.msl_altitudes" ;
    byte new_cal_trigger(calibration) ;
        new_cal_trigger:long_name = "Trigger of Calibration Change" ;
        new_cal_trigger:description = "reason for recalibration" ;
        new_cal_trigger:bit_0 = "radiosonde profile" ;
        new_cal_trigger:bit_1 = "i2 scan" ;
        new_cal_trigger:bit_2 = "geometry" ;
        new_cal_trigger:dpl_py_binding = "dne" ;
    short new_cal_offset(calibration) ;
        new_cal_offset:long_name = "Record Dimension equivalent Offset" ;
        new_cal_offset:min_value = 0 ;
        new_cal_offset:dpl_py_binding = "dne" ;
    float top_alt_sounding(calibration) ;
        top_alt_sounding:long_name = "Sounding Maximum Altitude" ;
        top_alt_sounding:units = "meters" ;
        top_alt_sounding:dpl_py_binding = "sounding.top" ;
    float raob_temperature(time, altitude) ;
        raob_temperature:long_name = "Raob Temperature Profile" ;
        raob_temperature:description = "Temperature interpolated to requested altitude resolution" ;
        raob_temperature:units = "degrees Kelvin" ;
        raob_temperature:dpl_py_binding = "rs_inv.temps" ;
    float raob_pressure(time, altitude) ;
        raob_pressure:long_name = "Raob pressure Profile" ;
        raob_pressure:description = "Pressure interpolated to requested altitude resolution" ;
        raob_pressure:units = "hectopascals" ;
        raob_pressure:dpl_py_binding = "rs_inv.pressures" ;
    float temperature_profile(calibration, altitude) ;
        temperature_profile:long_name = "Raob Temperature Profile" ;
        temperature_profile:description = "Temperature interpolated to requested altitude resolution" ;
        temperature_profile:units = "degrees Kelvin" ;
        temperature_profile:dpl_py_binding = "sounding.temps" ;
    float pressure_profile(calibration, altitude) ;
        pressure_profile:long_name = "Raob pressure Profile" ;
        pressure_profile:description = "Pressure interpolated to requested altitude resolution" ;
        pressure_profile:units = "hectopascals" ;
        pressure_profile:dpl_py_binding = "sounding.pressures" ;
    float dewpoint_profile(calibration, altitude) ;
        dewpoint_profile:long_name = "Raob Dewpoint Temperature Profile" ;
        dewpoint_profile:description = "Dewpoint interpolated to requested altitude resolution" ;
        dewpoint_profile:units = "degrees Kelvin" ;
        dewpoint_profile:missing_value = 9.96920996838687e+36 ;
        dewpoint_profile:dpl_py_binding = "sounding.dew_points" ;
    float windspeed_profile(calibration, altitude) ;
        windspeed_profile:long_name = "Raob Wind Speed Profile" ;
        windspeed_profile:description = "Speeds interpolated to requested altitude resolution" ;
        windspeed_profile:units = "m/s" ;
        windspeed_profile:missing_value = 9.96920996838687e+36 ;
        windspeed_profile:dpl_py_binding = "sounding.wind_spd" ;
    float winddir_profile(calibration, altitude) ;
        winddir_profile:long_name = "Raob Wind Direction Profile" ;
        winddir_profile:description = "Directions interpolated to requested altitude resolution" ;
        winddir_profile:units = "degrees" ;
        winddir_profile:missing_value = 9.96920996838687e+36 ;
        winddir_profile:dpl_py_binding = "sounding.wind_dir" ;
    char calibration_version(calibration, githash) ;
        calibration_version:long_name = "Calibration Tables GIT Version" ;
        calibration_version:dpl_py_binding = "gitversion" ;
    char raob_station(calibration, sondenamelength) ;
        raob_station:long_name = "Radiosonde Station ID" ;
        raob_station:dpl_py_binding = "sounding.sounding_id" ;
    char i2_txt_header(calibration, i2header) ;
        i2_txt_header:long_name = "i2_scan_file_text_info" ;
        i2_txt_header:description = "Contains name of file used to compute calibration" ;
        i2_txt_header:dpl_py_binding = "dne" ;
    char geo_txt_header(calibration, geoheader) ;
        geo_txt_header:long_name = "geometric_correction_file_txt_header." ;
        geo_txt_header:dpl_py_binding = "dne" ;
    char ap_txt_header(calibration, apheader) ;
        ap_txt_header:long_name = "afterpulse_correction_file_txt_header." ;
        ap_txt_header:dpl_py_binding = "dne" ;
    double raob_time_offset(calibration) ;
        raob_time_offset:units = "seconds" ;
        raob_time_offset:long_name = "Radiosonde Launch time offset" ;
        raob_time_offset:description = "Time after base time in seconds" ;
        raob_time_offset:dpl_py_binding = "dne" ;
    short raob_time_vector(calibration) ;
        raob_time_vector:long_name = "Radiosonde Launch time vector" ;
        raob_time_vector:description = "Time in [year month day hour min sec ms us] format" ;
        raob_time_vector:dpl_py_binding = "dne" ;
    float Cmc(calibration, altitude) ;
        Cmc:long_name = "Molecular in Combined Calibration" ;
        Cmc:dpl_py_binding = "rs_Cxx.Cmc" ;
    float Cmm(calibration, altitude) ;
        Cmm:long_name = "Molecular in Molecular Calibration" ;
        Cmm:dpl_py_binding = "rs_Cxx.Cmm" ;
    float Cmm_i2a(calibration, altitude) ;
        Cmm_i2a:long_name = "Molecular i2a in Molecular i2a Calibration" ;
        Cmm_i2a:dpl_py_binding = "rs_Cxx.Cmm_i2a" ;
    float Cam(calibration) ;
        Cam:long_name = "Aerosol in Molecular Calibration" ;
        Cam:dpl_py_binding = "rs_Cxx.Cam" ;
    float Cam_i2a(calibration) ;
        Cam_i2a:long_name = "Aerosol in Molecular i2a Calibration" ;
        Cam_i2a:dpl_py_binding = "rs_Cxx.Cam_i2a" ;
    float aeri_btemp_wavenumber(aeri_btemp_wavenumber) ;
        aeri_btemp_wavenumber:long_name = "Wave number" ;
        aeri_btemp_wavenumber:units = "cm^-1" ;
        aeri_btemp_wavenumber:missing_value = 9.96920996838687e+36 ;
        aeri_btemp_wavenumber:dpl_py_binding = "dne" ;
    float aeri_btemp(time, aeri_btemp_wavenumber) ;
        aeri_btemp:long_name = "AERI Brightness Temperature" ;
        aeri_btemp:units = "degK" ;
        aeri_btemp:missing_value = 9.96920996838687e+36 ;
        aeri_btemp:dpl_py_binding = "dne" ;
    float mwr_watervapor(time) ;
        mwr_watervapor:long_name = "MWR Water vapor along LOS path" ;
        mwr_watervapor:units = "cm" ;
        mwr_watervapor:missing_value = 9.96920996838687e+36 ;
        mwr_watervapor:dpl_py_binding = "dne" ;
    float mwr_liquidwater(time) ;
        mwr_liquidwater:long_name = "MWR Liquid water along LOS path" ;
        mwr_liquidwater:units = "g/m^2" ;
        mwr_liquidwater:missing_value = 9.96920996838687e+36 ;
        mwr_liquidwater:dpl_py_binding = "dne" ;
    float aeri_mean_rad_wavenumber_ch1(aeri_mean_rad_wavenumber_ch1) ;
        aeri_mean_rad_wavenumber_ch1:long_name = "Wave number" ;
        aeri_mean_rad_wavenumber_ch1:units = "cm^-1" ;
        aeri_mean_rad_wavenumber_ch1:missing_value = 9.96920996838687e+36 ;
        aeri_mean_rad_wavenumber_ch1:dpl_py_binding = "dne" ;
    float aeri1_mean_rad(time, aeri_mean_rad_wavenumber_ch1) ;
        aeri1_mean_rad:long_name = "Downwelling radiance interpolated to standard wavenumber scale Channel 1" ;
        aeri1_mean_rad:units = "mw/(m2 sr cm-1)" ;
        aeri1_mean_rad:missing_value = 9.96920996838687e+36 ;
        aeri1_mean_rad:dpl_py_binding = "dne" ;
    int aeri_qc(time) ;
        aeri_qc:long_name = "Aeri Quality" ;
        aeri_qc:bit_0 = "channel 1" ;
        aeri_qc:bit_1 = "channel 2" ;
        aeri_qc:missing_value = -1 ;
        aeri_qc:dpl_py_binding = "dne" ;
    float aeri_mean_rad_wavenumber_ch2(aeri_mean_rad_wavenumber_ch2) ;
        aeri_mean_rad_wavenumber_ch2:long_name = "Wave number" ;
        aeri_mean_rad_wavenumber_ch2:units = "cm^-1" ;
        aeri_mean_rad_wavenumber_ch2:missing_value = 9.96920996838687e+36 ;
        aeri_mean_rad_wavenumber_ch2:dpl_py_binding = "dne" ;
    float aeri2_mean_rad(time, aeri_mean_rad_wavenumber_ch2) ;
        aeri2_mean_rad:long_name = "Downwelling radiance interpolated to standard wavenumber scale Channel 2" ;
        aeri2_mean_rad:units = "mw/(m2 sr cm-1)" ;
        aeri2_mean_rad:missing_value = 9.96920996838687e+36 ;
        aeri2_mean_rad:dpl_py_binding = "dne" ;
    float aeri1_pca_mean_rad(time, aeri_mean_rad_wavenumber_ch1) ;
        aeri1_pca_mean_rad:long_name = "PCA Filtered Downwelling radiance interpolated to standard wavenumber scale Channel 1" ;
        aeri1_pca_mean_rad:units = "mw/(m2 sr cm-1)" ;
        aeri1_pca_mean_rad:missing_value = 9.96920996838687e+36 ;
        aeri1_pca_mean_rad:dpl_py_binding = "dne" ;
    float aeri2_pca_mean_rad(time, aeri_mean_rad_wavenumber_ch2) ;
        aeri2_pca_mean_rad:long_name = "PCA Filtered Downwelling radiance interpolated to standard wavenumber scale Channel 2" ;
        aeri2_pca_mean_rad:units = "mw/(m2 sr cm-1)" ;
        aeri2_pca_mean_rad:missing_value = 9.96920996838687e+36 ;
        aeri2_pca_mean_rad:dpl_py_binding = "dne" ;
    float beta_m(calibration, altitude) ;
        beta_m:long_name = "Raob molecular (Rayleigh) scattering cross section per unit volume" ;
        beta_m:units = "1/meter" ;
        beta_m:plot_scale = "logarithmic" ;
        beta_m:dpl_py_binding = "rs_Cxx.beta_r" ;
    float beta_m_1064(calibration, altitude) ;
        beta_m_1064:long_name = "Raob molecular (Rayleigh) 1064nm scattering cross section per unit volume" ;
        beta_m_1064:units = "1/meter" ;
        beta_m_1064:plot_scale = "logarithmic" ;
        beta_m_1064:dpl_py_binding = "rs_Cxx.beta_r_1064" ;
    float transmitted_energy(time) ;
        transmitted_energy:long_name = "Transmitted Energy" ;
        transmitted_energy:units = "Joules" ;
        transmitted_energy:missing_value = 9.96920996838687e+36 ;
        transmitted_energy:dpl_py_binding = "rs_mean.transmitted_energy" ;
    float transmitted_1064_energy(time) ;
        transmitted_1064_energy:long_name = "Transmitted 1064nm Energy" ;
        transmitted_1064_energy:units = "Joules" ;
        transmitted_1064_energy:missing_value = 9.96920996838687e+36 ;
        transmitted_1064_energy:dpl_py_binding = "rs_mean.transmitted_1064_energy" ;
    float piezovoltage(time) ;
        piezovoltage:long_name = "piezovoltage" ;
        piezovoltage:units = "Volts" ;
        piezovoltage:missing_value = 9.96920996838687e+36 ;
        piezovoltage:dpl_py_binding = "dne" ;
    int num_seeded_shots(time) ;
        num_seeded_shots:long_name = "Number of Seeded Shots" ;
        num_seeded_shots:missing_value = -1 ;
        num_seeded_shots:dpl_py_binding = "rs_mean.seeded_shots" ;
    int num_shots(time) ;
        num_shots:long_name = "Number of Shots" ;
        num_shots:missing_value = -1 ;
        num_shots:dpl_py_binding = "rs_mean.shot_count" ;
    float seed_quality(time) ;
        seed_quality:long_name = "Laser Seeding Quality" ;
        seed_quality:description = "The ratio of seeded shots to total shots. Only seeded shot data is stored and processed.  A low seed ratio can result in low noise resistance." ;
        seed_quality:missing_value = 9.96920996838687e+36 ;
        seed_quality:range = 0., 1. ;
        seed_quality:dpl_py_binding = "dne" ;
    float frequency_quality(time) ;
        frequency_quality:long_name = "Laser Frequency Quality" ;
        frequency_quality:description = "An ratio average of how good the frequency lock is per raw interval. A low value can result in poor separation of molecular and aerosol counts." ;
        frequency_quality:missing_value = 9.96920996838687e+36 ;
        frequency_quality:range = 0., 1. ;
        frequency_quality:dpl_py_binding = "dne" ;
    float lock_quality(time) ;
        lock_quality:long_name = "Laser Lock Quality" ;
        lock_quality:description = "A ratio of likely locked intervals (frequency_quality>=.5) to seeded intervals.  A low value can result in poor separation of molecular and aerosol counts." ;
        lock_quality:missing_value = 9.96920996838687e+36 ;
        lock_quality:range = 0., 1. ;
        lock_quality:dpl_py_binding = "dne" ;
    float mol_cal_pulse(time) ;
        mol_cal_pulse:long_name = "Molecular calibration pulse" ;
        mol_cal_pulse:description = "Sum of photon counts in the molecular channel due to light scattered with the telescope." ;
        mol_cal_pulse:units = "counts" ;
        mol_cal_pulse:missing_value = 9.96920996838687e+36 ;
        mol_cal_pulse:dpl_py_binding = "rs_mean.molecular_cal_pulse" ;
    float comb_hi_cal_pulse(time) ;
        comb_hi_cal_pulse:long_name = "Combined Hi calibration pulse" ;
        comb_hi_cal_pulse:description = "Sum of photon counts in the molecular channel due to light scattered with the telescope." ;
        comb_hi_cal_pulse:units = "counts" ;
        comb_hi_cal_pulse:missing_value = 9.96920996838687e+36 ;
        comb_hi_cal_pulse:dpl_py_binding = "rs_mean.combined_hi_cal_pulse" ;
    float comb_1064_cal_pulse(time) ;
        comb_1064_cal_pulse:long_name = "Combined 1064nm calibration pulse" ;
        comb_1064_cal_pulse:description = "Sum of photon counts in the molecular channel due to light scattered with the telescope." ;
        comb_1064_cal_pulse:units = "counts" ;
        comb_1064_cal_pulse:missing_value = 9.96920996838687e+36 ;
        comb_1064_cal_pulse:dpl_py_binding = "rs_mean.combined_1064_cal_pulse" ;
    int mol_norm_idx ;
        mol_norm_idx:dpl_py_binding = "rs_inv.mol_norm_index" ;
    float profile_num_seeded_shots(profile_time) ;
        profile_num_seeded_shots:long_name = "Profile Seeded shots" ;
        profile_num_seeded_shots:description = "Profile Seeded Shots" ;
        profile_num_seeded_shots:units = "shots" ;
        profile_num_seeded_shots:missing_value = 9.96920996838687e+36 ;
        profile_num_seeded_shots:dpl_py_binding = "profiles.seeded_shots" ;
    float profile_c_pol_dark_count(profile_time) ;
        profile_c_pol_dark_count:long_name = "Cross Polarization Dark Count FIXME dark counts need alt" ;
        profile_c_pol_dark_count:description = "Counts/bin at output resolution" ;
        profile_c_pol_dark_count:units = "counts" ;
        profile_c_pol_dark_count:missing_value = 9.96920996838687e+36 ;
        profile_c_pol_dark_count:dpl_py_binding = "profiles.c_pol_dark_counts" ;
    float profile_combined_1064_dark_count(profile_time) ;
        profile_combined_1064_dark_count:long_name = "Combined 1064nm Dark Count FIXME dark counts need alt" ;
        profile_combined_1064_dark_count:description = "Counts/bin at output resolution" ;
        profile_combined_1064_dark_count:units = "counts" ;
        profile_combined_1064_dark_count:missing_value = 9.96920996838687e+36 ;
        profile_combined_1064_dark_count:dpl_py_binding = "profiles.combined_1064_dark_counts" ;
    float profile_mol_dark_count(profile_time) ;
        profile_mol_dark_count:long_name = "Molecular Dark Count" ;
        profile_mol_dark_count:description = "Counts/bin at output resolution" ;
        profile_mol_dark_count:units = "counts" ;
        profile_mol_dark_count:missing_value = 9.96920996838687e+36 ;
        profile_mol_dark_count:dpl_py_binding = "profiles.mol_dark_counts" ;
    float profile_combined_dark_count_lo(profile_time) ;
        profile_combined_dark_count_lo:long_name = "Low Gain Combined Dark Count" ;
        profile_combined_dark_count_lo:description = "Counts/bin at output resolution" ;
        profile_combined_dark_count_lo:units = "counts" ;
        profile_combined_dark_count_lo:missing_value = 9.96920996838687e+36 ;
        profile_combined_dark_count_lo:dpl_py_binding = "profiles.c_lo_dark_counts" ;
    float profile_combined_dark_count_hi(profile_time) ;
        profile_combined_dark_count_hi:long_name = "High Gain Combined Dark Count" ;
        profile_combined_dark_count_hi:description = "Counts/bin at output resolution" ;
        profile_combined_dark_count_hi:units = "counts" ;
        profile_combined_dark_count_hi:missing_value = 9.96920996838687e+36 ;
        profile_combined_dark_count_hi:dpl_py_binding = "profiles.c_hi_dark_counts" ;
    float profile_mol_wfov_dark_count(profile_time) ;
        profile_mol_wfov_dark_count:long_name = "Molecular WFOV Dark Count" ;
        profile_mol_wfov_dark_count:description = "Counts/bin at output resolution" ;
        profile_mol_wfov_dark_count:units = "counts" ;
        profile_mol_wfov_dark_count:missing_value = 9.96920996838687e+36 ;
        profile_mol_wfov_dark_count:dpl_py_binding = "profiles.m_wfov_dark_counts" ;
    float profile_combined_wfov_dark_count(profile_time) ;
        profile_combined_wfov_dark_count:long_name = "Combined WFOV Dark Count" ;
        profile_combined_wfov_dark_count:description = "Counts/bin at output resolution" ;
        profile_combined_wfov_dark_count:units = "counts" ;
        profile_combined_wfov_dark_count:missing_value = 9.96920996838687e+36 ;
        profile_combined_wfov_dark_count:dpl_py_binding = "profiles.c_wfov_dark_counts" ;
    float profile_mol_i2a_dark_count(profile_time) ;
        profile_mol_i2a_dark_count:long_name = "Molecular I2A Dark Count" ;
        profile_mol_i2a_dark_count:description = "Counts/bin at output resolution" ;
        profile_mol_i2a_dark_count:units = "counts" ;
        profile_mol_i2a_dark_count:missing_value = 9.96920996838687e+36 ;
        profile_mol_i2a_dark_count:dpl_py_binding = "profiles.mol_i2a_dark_counts" ;
    float c_pol_dark_count(time) ;
        c_pol_dark_count:long_name = "Cross Polarization Dark Count FIXME dark counts need alt" ;
        c_pol_dark_count:description = "Counts/bin at output resolution" ;
        c_pol_dark_count:units = "counts" ;
        c_pol_dark_count:missing_value = 9.96920996838687e+36 ;
        c_pol_dark_count:dpl_py_binding = "rs_mean.c_pol_dark_counts" ;
    float mol_dark_count(time) ;
        mol_dark_count:long_name = "Molecular Dark Count" ;
        mol_dark_count:description = "Counts/bin at output resolution" ;
        mol_dark_count:units = "counts" ;
        mol_dark_count:missing_value = 9.96920996838687e+36 ;
        mol_dark_count:dpl_py_binding = "rs_mean.mol_dark_counts" ;
    float combined_dark_count_lo(time) ;
        combined_dark_count_lo:long_name = "Low Gain Combined Dark Count" ;
        combined_dark_count_lo:description = "Counts/bin at output resolution" ;
        combined_dark_count_lo:units = "counts" ;
        combined_dark_count_lo:missing_value = 9.96920996838687e+36 ;
        combined_dark_count_lo:dpl_py_binding = "rs_mean.c_lo_dark_counts" ;
    float combined_dark_count_1064(time) ;
        combined_dark_count_1064:long_name = "1064nm Combined Dark Count" ;
        combined_dark_count_1064:description = "Counts/bin at output resolution" ;
        combined_dark_count_1064:units = "counts" ;
        combined_dark_count_1064:missing_value = 9.96920996838687e+36 ;
        combined_dark_count_1064:dpl_py_binding = "rs_mean.combined_1064_dark_counts" ;
    float combined_dark_count_hi(time) ;
        combined_dark_count_hi:long_name = "High Gain Combined Dark Count" ;
        combined_dark_count_hi:description = "Counts/bin at output resolution" ;
        combined_dark_count_hi:units = "counts" ;
        combined_dark_count_hi:missing_value = 9.96920996838687e+36 ;
        combined_dark_count_hi:dpl_py_binding = "rs_mean.c_hi_dark_counts" ;
    float mol_wfov_dark_count(time) ;
        mol_wfov_dark_count:long_name = "Molecular WFOV Dark Count" ;
        mol_wfov_dark_count:description = "Counts/bin at output resolution" ;
        mol_wfov_dark_count:units = "counts" ;
        mol_wfov_dark_count:missing_value = 9.96920996838687e+36 ;
        mol_wfov_dark_count:dpl_py_binding = "rs_mean.m_wfov_dark_counts" ;
    float combined_wfov_dark_count(time) ;
        combined_wfov_dark_count:long_name = "Combined WFOV Dark Count" ;
        combined_wfov_dark_count:description = "Counts/bin at output resolution" ;
        combined_wfov_dark_count:units = "counts" ;
        combined_wfov_dark_count:missing_value = 9.96920996838687e+36 ;
        combined_wfov_dark_count:dpl_py_binding = "rs_mean.c_wfov_dark_counts" ;
    float mol_i2a_dark_count(time) ;
        mol_i2a_dark_count:long_name = "Molecular I2A Dark Count" ;
        mol_i2a_dark_count:description = "Counts/bin at output resolution" ;
        mol_i2a_dark_count:units = "counts" ;
        mol_i2a_dark_count:missing_value = 9.96920996838687e+36 ;
        mol_i2a_dark_count:dpl_py_binding = "rs_mean.mol_i2a_dark_counts" ;
    float combined_gain(calibration) ;
        combined_gain:long_name = "Combined Gain Factor" ;
        combined_gain:description = "Low Gain level * Factor ~ High Gain level" ;
        combined_gain:dpl_py_binding = "rs_constants.hi_to_low_combined_channel_gain_ratio" ;
    float combined_merge_threshhold(calibration) ;
        combined_merge_threshhold:long_name = "Combined Merge Threshhold" ;
        combined_merge_threshhold:dpl_py_binding = "rs_constants.combined_channel_merge_threshhold" ;
    float polarization_cross_talk(calibration) ;
        polarization_cross_talk:long_name = "Polarization Cross Talk" ;
        polarization_cross_talk:dpl_py_binding = "rs_constants.polarization_cross_talk" ;
    float wfov_to_combined_gain_ratio(calibration) ;
        wfov_to_combined_gain_ratio:long_name = "WFOV to Combined Gain" ;
        wfov_to_combined_gain_ratio:dpl_py_binding = "rs_constants.wfov_to_combined_gain_ratio" ;
    float combined_to_cross_pol_gain_ratio(calibration) ;
        combined_to_cross_pol_gain_ratio:long_name = "Combined to Cross Pol Gain" ;
        combined_to_cross_pol_gain_ratio:dpl_py_binding = "rs_constants.combined_to_cross_pol_gain_ratio" ;
    float molecular_to_wfov_gain_ratio(calibration) ;
        molecular_to_wfov_gain_ratio:long_name = "Molecular to WFOV Gain" ;
        molecular_to_wfov_gain_ratio:dpl_py_binding = "rs_constants.molecular_to_wfov_gain_ratio" ;
    float geo_cor(calibration, bin_range) ;
        geo_cor:long_name = "Overlap correction" ;
        geo_cor:description = "Geometric overlap correction in raw range bins" ;
        geo_cor:units = " " ;
        geo_cor:missing_value = 9.96920996838687e+36 ;
        geo_cor:plot_scale = "logarithmic" ;
        geo_cor:dpl_py_binding = "geo_corr" ;
    int od_norm_index ;
        od_norm_index:long_name = "Optical depth normalization index FIXME shouldn't be needed" ;
        od_norm_index:dpl_py_binding = "rs_inv.od_norm_index" ;
    int mol_ref_aod(time) ;
        mol_ref_aod:long_name = "optical depth below molecular reference altitude" ;
        mol_ref_aod:units = " " ;
        mol_ref_aod:description = "Estimated unmeasured optical depth below reference altitude--from linear extrapolation of extinction" ;
        mol_ref_aod:dpl_py_binding = "rs_inv.mol_ref_aod" ;
    float od(time, altitude) ;
        od:long_name = "Aerosol + Molecular Optical Depth" ;
        od:units = " " ;
        od:missing_value = 9.96920996838687e+36 ;
        od:insufficient_data = 9.96920996838687e+36 ;
        od:plot_scale = "logarithmic" ;
        od:dpl_py_binding = "rs_inv.optical_depth" ;
    float profile_std_beta_a_backscat(profile_time, altitude) ;
        profile_std_beta_a_backscat:long_name = "Std dev of backscat cross section (photon counting)" ;
        profile_std_beta_a_backscat:units = "1/(m sr)" ;
        profile_std_beta_a_backscat:missing_value = 9.96920996838687e+36 ;
        profile_std_beta_a_backscat:plot_scale = "logarithmic" ;
        profile_std_beta_a_backscat:dpl_py_binding = "profiles.inv.std_beta_a_backscat" ;
    float profile_od(profile_time,altitude) ;
        profile_od:long_name = "Aerosol + Molecular Optical Depth" ;
        profile_od:units = " " ;
        profile_od:missing_value = 9.96920996838687e+36 ;
        profile_od:insufficient_data = 9.96920996838687e+36 ;
        profile_od:plot_scale = "logarithmic" ;
        profile_od:dpl_py_binding = "profiles.inv.optical_depth" ;
    float od_aerosol(time, altitude) ;
        od_aerosol:long_name = "Aerosol Optical Depth" ;
        od_aerosol:units = " " ;
        od_aerosol:missing_value = 9.96920996838687e+36 ;
        od_aerosol:insufficient_data = 9.96920996838687e+36 ;
        od_aerosol:plot_scale = "logarithmic" ;
        od_aerosol:dpl_py_binding = "rs_inv.optical_depth_aerosol" ;
    float profile_od_aerosol(profile_time,altitude) ;
        profile_od_aerosol:long_name = "Aerosol Optical Depth" ;
        profile_od_aerosol:units = " " ;
        profile_od_aerosol:missing_value = 9.96920996838687e+36 ;
        profile_od_aerosol:insufficient_data = 9.96920996838687e+36 ;
        profile_od_aerosol:plot_scale = "logarithmic" ;
        profile_od_aerosol:dpl_py_binding = "profiles.inv.optical_depth_aerosol" ;
    float profile_extinction(profile_time,altitude) ;
        profile_extinction:long_name = "Aerosol + Molecular Extinction Profile" ;
        profile_extinction:units = " " ;
        profile_extinction:missing_value = 9.96920996838687e+36 ;
        profile_extinction:insufficient_data = 9.96920996838687e+36 ;
        profile_extinction:plot_scale = "logarithmic" ;
        profile_extinction:dpl_py_binding = "profiles.inv.extinction" ;
    float extinction(time,altitude) ;
        extinction:long_name = "Aerosol + Molecular Extinction" ;
        extinction:units = " " ;
        extinction:missing_value = 9.96920996838687e+36 ;
        extinction:insufficient_data = 9.96920996838687e+36 ;
        extinction:plot_scale = "logarithmic" ;
        extinction:dpl_py_binding = "rs_inv.extinction" ;
    float profile_extinction_aerosol(profile_time,altitude) ;
        profile_extinction_aerosol:long_name = "Aerosol Extinction Profile" ;
        profile_extinction_aerosol:units = " " ;
        profile_extinction_aerosol:missing_value = 9.96920996838687e+36 ;
        profile_extinction_aerosol:insufficient_data = 9.96920996838687e+36 ;
        profile_extinction_aerosol:plot_scale = "logarithmic" ;
        profile_extinction_aerosol:dpl_py_binding = "profiles.inv.extinction_aerosol" ;
    float extinction_aerosol(time,altitude) ;
        extinction_aerosol:long_name = "Aerosol Extinction" ;
        extinction_aerosol:units = " " ;
        extinction_aerosol:missing_value = 9.96920996838687e+36 ;
        extinction_aerosol:insufficient_data = 9.96920996838687e+36 ;
        extinction_aerosol:plot_scale = "logarithmic" ;
        extinction_aerosol:dpl_py_binding = "rs_inv.extinction_aerosol" ;
    float radar_backscattercrosssection(time, altitude) ;
        radar_backscattercrosssection:long_name = "Radar Backscatter Cross Section" ;
        radar_backscattercrosssection:units = "1/(m sr)" ;
        radar_backscattercrosssection:missing_value = 9.96920996838687e+36 ;
        radar_backscattercrosssection:dpl_py_binding = "rs_mmcr.Backscatter" ;
    float radar_reflectivity(time, altitude) ;
        radar_reflectivity:long_name = "Radar Reflectivity" ;
        radar_reflectivity:units = "dBz" ;
        radar_reflectivity:missing_value = 9.96920996838687e+36 ;
        radar_reflectivity:dpl_py_binding = "rs_mmcr.Reflectivity" ;
    float radar_spectralwidth(time, altitude) ;
        radar_spectralwidth:long_name = "Radar Spectral Width" ;
        radar_spectralwidth:units = "m/s" ;
        radar_spectralwidth:missing_value = 9.96920996838687e+36 ;
        radar_spectralwidth:dpl_py_binding = "rs_mmcr.SpectralWidth" ;
    float radar_dopplervelocity(time, altitude) ;
        radar_dopplervelocity:long_name = "Radar doppler Velocity" ;
        radar_dopplervelocity:units = "m/s" ;
        radar_dopplervelocity:missing_value = 9.96920996838687e+36 ;
        radar_dopplervelocity:dpl_py_binding = "rs_mmcr.MeanDopplerVelocity" ;
    float effective_diameter_prime(time, altitude) ;
        effective_diameter_prime:long_name = "lidar/radar effective particle diameter prime measurement" ;
        effective_diameter_prime:units = "m" ;
        effective_diameter_prime:description = "Effective diameter directly from the ratio of Lidar Backscatter and Radar Reflectivity; (<volume^2>/<area>)^.25, see Donovan JGR Nov 2001" ;
        effective_diameter_prime:missing_value = 9.96920996838687e+36 ;
        effective_diameter_prime:dpl_py_binding = "rs_spheroid_particle.effective_diameter_prime" ;
    float effective_diameter(time, altitude) ;
        effective_diameter:long_name = "Effective particle diameter" ;
        effective_diameter:units = "m" ;
        effective_diameter:description = "Effective particle diameter derived from ratio of Lidar Backscatter and Radar Reflectivity; assuming a gamma size distribution using assumptions from particle processing parameters" ;
        effective_diameter:missing_value = 9.96920996838687e+36 ;
        effective_diameter:dpl_py_binding = "rs_spheroid_particle.effective_diameter" ;
    float num_particles(time, altitude) ;
        num_particles:long_name = "Number density of particles" ;
        num_particles:units = "1/liter" ;
        num_particles:description = "Number of particles per liter derived from ratio of lidar backscatter and radar reflectivity; assuming a gamma size distribution" ;
        num_particles:missing_value = 9.96920996838687e+36 ;
        num_particles:dpl_py_binding = "rs_spheroid_particle.num_particles" ;
    float mean_diameter(time, altitude) ;
        mean_diameter:long_name = "Mean diameter of particles" ;
        mean_diameter:units = "m" ;
        mean_diameter:description = "Mean diameter of particles derived from the effective diameter and the gamma size distribution" ;
        mean_diameter:missing_value = 9.96920996838687e+36 ;
        mean_diameter:dpl_py_binding = "rs_spheroid_particle.mean_diameter" ;
    float LWC(time, altitude) ;
        LWC:long_name = "Liquid water content" ;
        LWC:units = "kg/m^3" ;
        LWC:description = "Liquid water content derived from ratio of lidar backscatter and radar reflectivity; assuming a gamma size distribution" ;
        LWC:missing_value = 9.96920996838687e+36 ;
        LWC:dpl_py_binding = "rs_spheroid_particle.LWC" ;
    float precip_rate(time, altitude) ;
        precip_rate:long_name = "HSRL-Radar Precipitation Rate" ;
        precip_rate:units = "m/s" ;
        precip_rate:description = "precipitation accumulation rate from combined hsrl radar retrieval" ;
        precip_rate:missing_value = 9.96920996838687e+36 ;
        precip_rate:dpl_py_binding = "rs_spheroid_particle.hsrl_radar_precip_rate" ;
    float fall_velocity(time, altitude) ;
        fall_velocity:long_name = "radar-weighted fall velocity" ;
        fall_velocity:units = "m/s" ;
        fall_velocity:description = "modeled fall velocity weighted by radar cross section" ;
        fall_velocity:missing_value = 9.96920996838687e+36 ;
        fall_velocity:dpl_py_binding = "rs_spheroid_particle.rw_fall_velocity" ;
    float model_spectral_width(time, altitude) ;
        model_spectral_width:long_name = "Modeled Radar Spectral Width" ;
        model_spectral_width:units = "m/s" ;
        model_spectral_width:description = "radar spectral width modeled from derived hsrl_radar particle size retrieval" ;
        model_spectral_width:missing_value = 9.96920996838687e+36 ;
        model_spectral_width:dpl_py_binding = "rs_spheroid_particle.model_spectral_width" ;
    float beta_a(time, altitude) ;
        beta_a:long_name = "Particulate extinction cross section per unit volume" ;
        beta_a:units = "1/m" ;
        beta_a:missing_value = 9.96920996838687e+36 ;
        beta_a:plot_scale = "logarithmic" ;
        beta_a:dpl_py_binding = "rs_inv.beta_a" ;
    float integrated_backscat(time, altitude) ;
        integrated_backscat:long_name = "Range-integrated backscatter cross section" ;
        integrated_backscat:units = "1/sr" ;
        integrated_backscat:missing_value = 9.96920996838687e+36 ;
        integrated_backscat:plot_scale = "logarithmic" ;
        integrated_backscat:dpl_py_binding = "rs_inv.integrated_backscatter" ;
    float atten_beta_a_backscat(time, altitude) ;
        atten_beta_a_backscat:long_name = "Attenuated Molecular return" ;
        atten_beta_a_backscat:units = "1/(m sr)" ;
        atten_beta_a_backscat:missing_value = 9.96920996838687e+36 ;
        atten_beta_a_backscat:plot_scale = "logarithmic" ;
        atten_beta_a_backscat:dpl_py_binding = "rs_inv.atten_beta_a_backscat" ;
    float atten_beta_a_1064_backscat(time, altitude) ;
        atten_beta_a_1064_backscat:long_name = "Attenuated 1064nm Molecular return" ;
        atten_beta_a_1064_backscat:units = "1/(m sr)" ;
        atten_beta_a_1064_backscat:missing_value = 9.96920996838687e+36 ;
        atten_beta_a_1064_backscat:plot_scale = "logarithmic" ;
        atten_beta_a_1064_backscat:dpl_py_binding = "rs_inv.attenuated_1064_backscatter" ;
    float profile_atten_beta_a_backscat(altitude) ;
        profile_atten_beta_a_backscat:long_name = "Attenuated Molecular Profile" ;
        profile_atten_beta_a_backscat:units = "1/(m sr)" ;
        profile_atten_beta_a_backscat:missing_value = 9.96920996838687e+36 ;
        profile_atten_beta_a_backscat:plot_scale = "logarithmic" ;
        profile_atten_beta_a_backscat:dpl_py_binding = "profiles.inv.atten_beta_a_backscat" ;
    float circular_depol(time, altitude) ;
        circular_depol:long_name = "Circular depolarization ratio for particulate" ;
        circular_depol:description = "left circular return divided by right circular return" ;
        circular_depol:units = "%" ;
        circular_depol:missing_value = 9.96920996838687e+36 ;
        circular_depol:plot_scale = "logarithmic" ;
        circular_depol:dpl_py_binding = "rs_inv.circular_depol" ;
    float linear_depol_i2a(time, altitude) ;
        linear_depol_i2a:long_name = "Linear depolarization i2a ratio for particulate" ;
        linear_depol_i2a:description = "Perpendicular / parallel_i2a polarization" ;
        linear_depol_i2a:units = "%" ;
        linear_depol_i2a:missing_value = 9.96920996838687e+36 ;
        linear_depol_i2a:plot_scale = "logarithmic" ;
        linear_depol_i2a:dpl_py_binding = "rs_inv.linear_depol_i2a" ;
    float linear_depol(time, altitude) ;
        linear_depol:long_name = "Linear depolarization ratio for particulate" ;
        linear_depol:description = "Perpendicular / parallel polarization" ;
        linear_depol:units = "%" ;
        linear_depol:missing_value = 9.96920996838687e+36 ;
        linear_depol:plot_scale = "logarithmic" ;
        linear_depol:dpl_py_binding = "rs_inv.linear_depol" ;
    float profile_circular_depol(profile_time,altitude) ;
        profile_circular_depol:long_name = "Circular depolarization ratio profile for particulate" ;
        profile_circular_depol:description = "left circular return divided by right circular return" ;
        profile_circular_depol:units = "%" ;
        profile_circular_depol:missing_value = 9.96920996838687e+36 ;
        profile_circular_depol:plot_scale = "logarithmic" ;
        profile_circular_depol:dpl_py_binding = "profiles.inv.circular_depol" ;
    float profile_linear_depol_i2a(profile_time,altitude) ;
        profile_linear_depol_i2a:long_name = "Linear depolarization i2a ratio profile for particulate" ;
        profile_linear_depol_i2a:description = "Perpendicular / parallel_i2a polarization" ;
        profile_linear_depol_i2a:units = "%" ;
        profile_linear_depol_i2a:missing_value = 9.96920996838687e+36 ;
        profile_linear_depol_i2a:plot_scale = "logarithmic" ;
        profile_linear_depol_i2a:dpl_py_binding = "profiles.inv.linear_depol_i2a" ;
    float profile_linear_depol(profile_time,altitude) ;
        profile_linear_depol:long_name = "Linear depolarization ratio profile for particulate" ;
        profile_linear_depol:description = "Perpendicular / parallel polarization" ;
        profile_linear_depol:units = "%" ;
        profile_linear_depol:missing_value = 9.96920996838687e+36 ;
        profile_linear_depol:plot_scale = "logarithmic" ;
        profile_linear_depol:dpl_py_binding = "profiles.inv.linear_depol" ;
    int molecular_wfov_counts(raw_time, bin_range) ;
        molecular_wfov_counts:long_name = "Molecular WFOV Photon Counts" ;
        molecular_wfov_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
        molecular_wfov_counts:units = "counts" ;
        molecular_wfov_counts:missing_value = -1 ;
        molecular_wfov_counts:plot_scale = "logarithmic" ;
        molecular_wfov_counts:dpl_py_binding = "rs_raw.molecular_wfov_counts" ;
    float profile_molecular_wfov_counts(profile_time,altitude) ;
        profile_molecular_wfov_counts:long_name = "Molecular WFOV Photon Counts profile" ;
        profile_molecular_wfov_counts:description = "Raw counts profile with pileup, afterpulse, and darkcount corrections applied" ;
        profile_molecular_wfov_counts:units = "counts" ;
        profile_molecular_wfov_counts:missing_value = -1 ;
        profile_molecular_wfov_counts:plot_scale = "logarithmic" ;
        profile_molecular_wfov_counts:dpl_py_binding = "profiles.molecular_wfov_counts" ;
    float profile_raw_molecular_wfov_counts(profile_time,bin_range) ;
        profile_raw_molecular_wfov_counts:long_name = "Raw Molecular WFOV Photon Counts profile" ;
        profile_raw_molecular_wfov_counts:description = "Raw counts profile with pileup" ;
        profile_raw_molecular_wfov_counts:units = "counts" ;
        profile_raw_molecular_wfov_counts:missing_value = -1 ;
        profile_raw_molecular_wfov_counts:plot_scale = "logarithmic" ;
        profile_raw_molecular_wfov_counts:dpl_py_binding = "profiles.raw_molecular_wfov_counts" ;
    int molecular_i2a_counts(raw_time, bin_range) ;
        molecular_i2a_counts:long_name = "Molecular Argon Photon Counts" ;
        molecular_i2a_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
        molecular_i2a_counts:units = "counts" ;
        molecular_i2a_counts:missing_value = -1 ;
        molecular_i2a_counts:plot_scale = "logarithmic" ;
        molecular_i2a_counts:dpl_py_binding = "rs_raw.molecular_i2a_counts" ;
    float profile_molecular_i2a_counts(profile_time,altitude) ;
        profile_molecular_i2a_counts:long_name = "Molecular Argon Photon Counts profile" ;
        profile_molecular_i2a_counts:description = "Raw counts profile with pileup, afterpulse, and darkcount corrections applied" ;
        profile_molecular_i2a_counts:units = "counts" ;
        profile_molecular_i2a_counts:missing_value = -1 ;
        profile_molecular_i2a_counts:plot_scale = "logarithmic" ;
        profile_molecular_i2a_counts:dpl_py_binding = "profiles.molecular_i2a_counts" ;
    float profile_raw_molecular_i2a_counts(profile_time,bin_range) ;
        profile_raw_molecular_i2a_counts:long_name = "Raw Molecular Argon Photon Counts profile" ;
        profile_raw_molecular_i2a_counts:description = "Raw counts profile with pileup" ;
        profile_raw_molecular_i2a_counts:units = "counts" ;
        profile_raw_molecular_i2a_counts:missing_value = -1 ;
        profile_raw_molecular_i2a_counts:plot_scale = "logarithmic" ;
        profile_raw_molecular_i2a_counts:dpl_py_binding = "profiles.raw_molecular_i2a_counts" ;
    int molecular_counts(raw_time, bin_range) ;
        molecular_counts:long_name = "Molecular Photon Counts" ;
        molecular_counts:description = "Raw counts profile with pileup correction applied" ;
        molecular_counts:units = "counts" ;
        molecular_counts:missing_value = -1 ;
        molecular_counts:plot_scale = "logarithmic" ;
        molecular_counts:dpl_py_binding = "rs_raw.molecular_counts" ;
    float profile_molecular_counts(profile_time,altitude) ;
        profile_molecular_counts:long_name = "Molecular Photon Counts profile" ;
        profile_molecular_counts:description = "Raw counts profile with pileup, afterpulse, and darkcount corrections applied" ;
        profile_molecular_counts:units = "counts" ;
        profile_molecular_counts:missing_value = -1 ;
        profile_molecular_counts:plot_scale = "logarithmic" ;
        profile_molecular_counts:dpl_py_binding = "profiles.molecular_counts" ;
    float profile_raw_molecular_counts(profile_time,bin_range) ;
        profile_raw_molecular_counts:long_name = "Raw Molecular Photon Counts profile" ;
        profile_raw_molecular_counts:description = "Raw counts profile with pileup applied" ;
        profile_raw_molecular_counts:units = "counts" ;
        profile_raw_molecular_counts:missing_value = -1 ;
        profile_raw_molecular_counts:plot_scale = "logarithmic" ;
        profile_raw_molecular_counts:dpl_py_binding = "profiles.raw_molecular_counts" ;
    int combined_counts_lo(raw_time, bin_range) ;
        combined_counts_lo:long_name = "Low Gain Combined Photon Counts" ;
        combined_counts_lo:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
        combined_counts_lo:units = "counts" ;
        combined_counts_lo:missing_value = -1 ;
        combined_counts_lo:plot_scale = "logarithmic" ;
        combined_counts_lo:dpl_py_binding = "rs_raw.combined_lo_counts" ;
    int combined_counts_hi(raw_time, bin_range) ;
        combined_counts_hi:long_name = "High Gain Combined Photon Counts" ;
        combined_counts_hi:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
        combined_counts_hi:units = "counts" ;
        combined_counts_hi:missing_value = -1 ;
        combined_counts_hi:plot_scale = "logarithmic" ;
        combined_counts_hi:dpl_py_binding = "rs_raw.combined_hi_counts" ;
    int combined_counts_1064(raw_time, bin_range) ;
        combined_counts_1064:long_name = "1064nm Combined Photon Counts" ;
        combined_counts_1064:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
        combined_counts_1064:units = "counts" ;
        combined_counts_1064:missing_value = -1 ;
        combined_counts_1064:plot_scale = "logarithmic" ;
        combined_counts_1064:dpl_py_binding = "rs_raw.combined_1064_counts" ;
    float profile_combined_counts_lo(profile_time,altitude) ;
        profile_combined_counts_lo:long_name = "Low Gain Combined Photon Counts profile" ;
        profile_combined_counts_lo:description = "Raw counts profile with pileup, afterpulse, and darkcount corrections applied" ;
        profile_combined_counts_lo:units = "counts" ;
        profile_combined_counts_lo:missing_value = -1 ;
        profile_combined_counts_lo:plot_scale = "logarithmic" ;
        profile_combined_counts_lo:dpl_py_binding = "profiles.combined_lo_counts" ;
    float profile_combined_counts_hi(profile_time,altitude) ;
        profile_combined_counts_hi:long_name = "High Gain Combined Photon Counts profile" ;
        profile_combined_counts_hi:description = "Raw counts profile with pileup, afterpulse, and darkcount corrections applied" ;
        profile_combined_counts_hi:units = "counts" ;
        profile_combined_counts_hi:missing_value = -1 ;
        profile_combined_counts_hi:plot_scale = "logarithmic" ;
        profile_combined_counts_hi:dpl_py_binding = "profiles.combined_hi_counts" ;
    float profile_combined_1064_counts(profile_time,altitude) ;
        profile_combined_1064_counts:long_name = "1064nm Combined Photon Counts profile" ;
        profile_combined_1064_counts:description = "Raw counts profile with pileup, afterpulse, and darkcount corrections applied" ;
        profile_combined_1064_counts:units = "counts" ;
        profile_combined_1064_counts:missing_value = -1 ;
        profile_combined_1064_counts:plot_scale = "logarithmic" ;
        profile_combined_1064_counts:dpl_py_binding = "profiles.combined_1064_counts" ;
    int cross_counts(raw_time, bin_range) ;
        cross_counts:long_name = "Cross Polarized Photon Counts" ;
        cross_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
        cross_counts:units = "counts" ;
        cross_counts:missing_value = -1 ;
        cross_counts:plot_scale = "logarithmic" ;
        cross_counts:dpl_py_binding = "rs_raw.cross_pol_counts" ;
    float profile_cross_counts(profile_time,altitude) ;
        profile_cross_counts:long_name = "Cross Polarized Photon Counts profile" ;
        profile_cross_counts:description = "Raw counts profile with pileup, afterpulse, and darkcount corrections applied" ;
        profile_cross_counts:units = "counts" ;
        profile_cross_counts:missing_value = -1 ;
        profile_cross_counts:plot_scale = "logarithmic" ;
        profile_cross_counts:dpl_py_binding = "profiles.cross_pol_counts" ;
    float beta_a_backscat_parallel(time, altitude) ;
        beta_a_backscat_parallel:long_name = "Particulate nondepolarized backscatter cross section per unit volume" ;
        beta_a_backscat_parallel:units = "1/(m sr)" ;
        beta_a_backscat_parallel:missing_value = 9.96920996838687e+36 ;
        beta_a_backscat_parallel:plot_scale = "logarithmic" ;
        beta_a_backscat_parallel:dpl_py_binding = "rs_inv.beta_a_backscat_par" ;
    float profile_beta_a_backscat_parallel(profile_time,altitude) ;
        profile_beta_a_backscat_parallel:long_name = "Particulate nondepolarized backscatter cross section profile" ;
        profile_beta_a_backscat_parallel:units = "1/(m sr)" ;
        profile_beta_a_backscat_parallel:missing_value = 9.96920996838687e+36 ;
        profile_beta_a_backscat_parallel:plot_scale = "logarithmic" ;
        profile_beta_a_backscat_parallel:dpl_py_binding = "profiles.inv.beta_a_backscat_par" ;
    float beta_a_backscat_perpendicular(time, altitude) ;
        beta_a_backscat_perpendicular:long_name = "Particulate depolarized backscatter cross section per unit volume" ;
        beta_a_backscat_perpendicular:units = "1/(m sr)" ;
        beta_a_backscat_perpendicular:missing_value = 9.96920996838687e+36 ;
        beta_a_backscat_perpendicular:plot_scale = "logarithmic" ;
        beta_a_backscat_perpendicular:dpl_py_binding = "rs_inv.beta_a_backscat_perp" ;
    float profile_beta_a_backscat_perpendicular(profile_time,altitude) ;
        profile_beta_a_backscat_perpendicular:long_name = "Particulate depolarized backscatter cross section profile" ;
        profile_beta_a_backscat_perpendicular:units = "1/(m sr)" ;
        profile_beta_a_backscat_perpendicular:missing_value = 9.96920996838687e+36 ;
        profile_beta_a_backscat_perpendicular:plot_scale = "logarithmic" ;
        profile_beta_a_backscat_perpendicular:dpl_py_binding = "profiles.inv.beta_a_backscat_perp" ;
    float beta_a_backscat(time, altitude) ;
        beta_a_backscat:long_name = "Particulate backscatter cross section per unit volume" ;
        beta_a_backscat:units = "1/(m sr)" ;
        beta_a_backscat:missing_value = 9.96920996838687e+36 ;
        beta_a_backscat:plot_scale = "logarithmic" ;
        beta_a_backscat:dpl_py_binding = "rs_inv.beta_a_backscat" ;
    float beta_a_1064_backscat(time, altitude) ;
        beta_a_1064_backscat:long_name = "Particulate 1064nm backscatter cross section per unit volume" ;
        beta_a_1064_backscat:units = "1/(m sr)" ;
        beta_a_1064_backscat:missing_value = 9.96920996838687e+36 ;
        beta_a_1064_backscat:plot_scale = "logarithmic" ;
        beta_a_1064_backscat:dpl_py_binding = "rs_inv.beta_a_1064_backscat" ;
    float profile_beta_a_backscat(profile_time,altitude) ;
        profile_beta_a_backscat:long_name = "Particulate backscatter cross section profile" ;
        profile_beta_a_backscat:units = "1/(m sr)" ;
        profile_beta_a_backscat:missing_value = 9.96920996838687e+36 ;
        profile_beta_a_backscat:plot_scale = "logarithmic" ;
        profile_beta_a_backscat:dpl_py_binding = "profiles.inv.beta_a_backscat" ;
    float profile_beta_a_1064_backscat(profile_time,altitude) ;
        profile_beta_a_1064_backscat:long_name = "Particulate 1064nm backscatter cross section profile" ;
        profile_beta_a_1064_backscat:units = "1/(m sr)" ;
        profile_beta_a_1064_backscat:missing_value = 9.96920996838687e+36 ;
        profile_beta_a_1064_backscat:plot_scale = "logarithmic" ;
        profile_beta_a_1064_backscat:dpl_py_binding = "profiles.inv.beta_a_1064_backscat" ;
    float Na_i2a(time, altitude) ;
        Na_i2a:long_name = "Inverted Aerosol Argon" ;
        Na_i2a:units = " " ;
        Na_i2a:dpl_py_binding = "rs_inv.Na_i2a" ;
    float Nm_i2a(time, altitude) ;
        Nm_i2a:long_name = "Inverted Molecular Argon" ;
        Nm_i2a:units = " " ;
        Nm_i2a:dpl_py_binding = "rs_inv.Nm_i2a" ;
    float Ncp_i2a(time, altitude) ;
        Ncp_i2a:long_name = "Inverted Cross Polarization Argon" ;
        Ncp_i2a:units = " " ;
        Ncp_i2a:dpl_py_binding = "rs_inv.Ncp_i2a" ;
    float Na(time, altitude) ;
        Na:long_name = "Inverted Aerosol" ;
        Na:units = " " ;
        Na:dpl_py_binding = "rs_inv.Na" ;
    float Nm(time, altitude) ;
        Nm:long_name = "Inverted Molecular" ;
        Nm:units = " " ;
        Nm:dpl_py_binding = "rs_inv.Nm" ;
    float Ncp(time, altitude) ;
        Ncp:long_name = "Inverted Cross Polarization" ;
        Ncp:units = " " ;
        Ncp:dpl_py_binding = "rs_inv.Ncp" ;
    float profile_Na(profile_time,altitude) ;
        profile_Na:long_name = "Inverted Aerosol Profile" ;
        profile_Na:units = " " ;
        profile_Na:dpl_py_binding = "profiles.inv.Na" ;
    float profile_Nm(profile_time,altitude) ;
        profile_Nm:long_name = "Inverted Molecular Profile" ;
        profile_Nm:units = " " ;
        profile_Nm:dpl_py_binding = "profiles.inv.Nm" ;
    float profile_Ncp(profile_time,altitude) ;
        profile_Ncp:long_name = "Inverted Cross Polarization Profile" ;
        profile_Ncp:units = " " ;
        profile_Ncp:dpl_py_binding = "profiles.inv.Ncp" ;
    float profile_Na_i2a(profile_time,altitude) ;
        profile_Na_i2a:long_name = "Inverted Aerosol Argon Profile" ;
        profile_Na_i2a:units = " " ;
        profile_Na_i2a:dpl_py_binding = "profiles.inv.Na_i2a" ;
    float profile_Nm_i2a(profile_time,altitude) ;
        profile_Nm_i2a:long_name = "Inverted Molecular Argon Profile" ;
        profile_Nm_i2a:units = " " ;
        profile_Nm_i2a:dpl_py_binding = "profiles.inv.Nm_i2a" ;
    float profile_Ncp_i2a(profile_time,altitude) ;
        profile_Ncp_i2a:long_name = "Inverted Cross Polarization Argon Profile" ;
        profile_Ncp_i2a:units = " " ;
        profile_Ncp_i2a:dpl_py_binding = "profiles.inv.Ncp_i2a" ;
    float temperature_profile_i2a(altitude) ;
        temperature_profile_i2a:long_name = "HSRL Iodine-Argon Temperature Profile" ;
        temperature_profile_i2a:description = "Temperature profile extracted from ratio of Argon-broadened and non-broadened molecular signals across entire time interval" ;
        temperature_profile_i2a:units = "degK" ;
        temperature_profile_i2a:dpl_py_binding = "profiles.i2a_temperatures" ;
    int qc_mask(time, altitude) ;
        qc_mask:long_name = "Quality Mask" ;
        qc_mask:description = "Quality mask bitfield.  Unused bits are always high" ;
        qc_mask:missing_value = 0 ;
        qc_mask:_Unsigned = "true" ;
        qc_mask:bit_0 = "complete_mask" ;
        qc_mask:bit_0_description = "data is good.  and of bits 1-9" ;
        qc_mask:bit_1 = "lidar_ok_mask" ;
        qc_mask:bit_1_description = "lidar data is present" ;
        qc_mask:bit_2 = "lock_quality_mask" ;
        qc_mask:bit_2_description = "laser is locked to iodine filter wavelength" ;
        qc_mask:bit_3 = "seed_quality_mask" ;
        qc_mask:bit_3_description = "laser wavelength is locked to seed laser" ;
        qc_mask:bit_4 = "mol_count_snr_mask" ;
        qc_mask:bit_4_description = "molecular signal/photon counting error in molecular signal is above specified threshhold" ;
        qc_mask:bit_5 = "backscat_snr_mask" ;
        qc_mask:bit_5_description = "backscatter cross-section/photon counting error in backscatter cross-section is above specified threshhold" ;
        qc_mask:bit_6 = "mol_lost_mask" ;
        qc_mask:bit_6_description = "number of molecular photon counts is above specified threshhold" ;
        qc_mask:bit_7 = "min_backscat_mask" ;
        qc_mask:bit_7_description = "lidar backscatter cross-section is above specified threshhold" ;
        qc_mask:bit_8 = "radar_backscat_mask" ;
        qc_mask:bit_8_description = "radar backscatter cross-section is above specified threshhold" ;
        qc_mask:bit_9 = "radar_ok_mask" ;
        qc_mask:bit_9_description = "radar data is present" ;
        qc_mask:bit_10 = "aeri_ok_mask" ;
        qc_mask:bit_10_description = "aeri data is present" ;
        qc_mask:bit_11 = "aeri_qc_mask" ;
        qc_mask:bit_11_description = "aeri data has passed a quality check" ;
        qc_mask:bit_12 = "cloud_mask" ;
        qc_mask:bit_12_description = "cloud encountered" ;
        qc_mask:dpl_py_binding = "rs_inv.qc_mask" ;
    float molecular_signal_to_noise(time, altitude) ;
        molecular_signal_to_noise:long_name = "Molecular Signal-to-Noise" ;
        molecular_signal_to_noise:description = "Molecular Signal-to-Noise computed from photon statistics" ;
        molecular_signal_to_noise:units = "" ;
        molecular_signal_to_noise:missing_value = 9.96920996838687e+36 ;
        molecular_signal_to_noise:plot_scale = "logarithmic" ;
        molecular_signal_to_noise:dpl_py_binding = "rs_inv.SN_mol" ;
    float molecular_i2a_signal_to_noise(time, altitude) ;
        molecular_i2a_signal_to_noise:long_name = "Molecular I2A Signal-to-Noise" ;
        molecular_i2a_signal_to_noise:description = "Molecular I2A Signal-to-Noise computed from photon statistics" ;
        molecular_i2a_signal_to_noise:units = "" ;
        molecular_i2a_signal_to_noise:missing_value = 9.96920996838687e+36 ;
        molecular_i2a_signal_to_noise:plot_scale = "logarithmic" ;
        molecular_i2a_signal_to_noise:dpl_py_binding = "rs_inv.SN_i2a_mol" ;
    float particulate_backscatter_signal_to_noise(time, altitude) ;
        particulate_backscatter_signal_to_noise:long_name = "Particulate Backscatter Signal-to-Noise" ;
        particulate_backscatter_signal_to_noise:description = "Particulate Backscatter Signal-to-Noise computed from photon statistics" ;
        particulate_backscatter_signal_to_noise:units = "" ;
        particulate_backscatter_signal_to_noise:missing_value = 9.96920996838687e+36 ;
        particulate_backscatter_signal_to_noise:plot_scale = "logarithmic" ;
        particulate_backscatter_signal_to_noise:dpl_py_binding = "rs_inv.SN_beta_a_backscat" ;
    float std_backscatter_ratio(time, altitude) ;
        std_backscatter_ratio:long_name = "Standard Deviation of Backscatter Ratio" ;
        std_backscatter_ratio:description = "Standard Deviation of Backscatter Ratio computed from photon statistics" ;
        std_backscatter_ratio:units = "" ;
        std_backscatter_ratio:missing_value = 9.96920996838687e+36 ;
        std_backscatter_ratio:plot_scale = "logarithmic" ;
        std_backscatter_ratio:dpl_py_binding = "rs_inv.SR_std" ;
    float std_beta_a_backscat(time, altitude) ;
        std_beta_a_backscat:long_name = "Std dev of backscat cross section (photon counting)" ;
        std_beta_a_backscat:units = "1/(m sr)" ;
        std_beta_a_backscat:missing_value = 9.96920996838687e+36 ;
        std_beta_a_backscat:plot_scale = "logarithmic" ;
        std_beta_a_backscat:dpl_py_binding = "rs_inv.std_beta_a_backscat" ;
    float mwr_frequency(mwr_frequency) ;
        mwr_frequency:long_name = "Frequency" ;
        mwr_frequency:units = "GHz" ;
        mwr_frequency:missing_value = 9.96920996838687e+36 ;
        mwr_frequency:dpl_py_binding = "dne" ;
    float mwr_btemp(time, mwr_frequency) ;
        mwr_btemp:long_name = "MWR Brightness Temperature" ;
        mwr_btemp:units = "degK" ;
        mwr_btemp:missing_value = 9.96920996838687e+36 ;
        mwr_btemp:dpl_py_binding = "dne" ;
    short hsrl_qa_BS(time, altitude) ;
        hsrl_qa_BS:long_name = "Quality Assurance Backscatter" ;
        hsrl_qa_BS:value_NC = 0 ;
        hsrl_qa_BS:value_Good = 1 ;
        hsrl_qa_BS:value_Bad = 2 ;
        hsrl_qa_BS:value_Caution = 3 ;
        hsrl_qa_BS:dpl_py_binding = "rs_inv.qa_flags.qa_BS" ;
    short hsrl_qa_dep(time, altitude) ;
        hsrl_qa_dep:long_name = "Quality Assurance Depolarization" ;
        hsrl_qa_dep:value_NC = 0 ;
        hsrl_qa_dep:value_Good = 1 ;
        hsrl_qa_dep:value_Bad = 2 ;
        hsrl_qa_dep:value_Caution = 3 ;
        hsrl_qa_dep:dpl_py_binding = "rs_inv.qa_flags.qa_dep" ;
    short hsrl_qa_Ext(time, altitude) ;
        hsrl_qa_Ext:long_name = "Quality Assurance Extinction" ;
        hsrl_qa_Ext:value_NC = 0 ;
        hsrl_qa_Ext:value_Good = 1 ;
        hsrl_qa_Ext:value_Bad = 2 ;
        hsrl_qa_Ext:value_Caution = 3 ;
        hsrl_qa_Ext:dpl_py_binding = "rs_inv.qa_flags.qa_Ext" ;
        
    float rlprof_asr(time, altitude) ;
        rlprof_asr:long_name = "Raman Aerosol Scattering Ratio" ;
        rlprof_asr:units = "unitless" ;
        rlprof_asr:dpl_py_binding = "rlprofaerosol.aerosol_backscatter_ratio" ;
    float rlprof_asr_error(time, altitude) ;
        rlprof_asr_error:long_name = "Uncertainty in calibrated aerosol scattering ratio" ;
        rlprof_asr_error:units = "unitless" ;
        rlprof_asr_error:dpl_py_binding = "rlprofaerosol.aerosol_backscatter_ratio_error" ;
    float rlprof_beta(time, altitude) ;
        rlprof_beta:long_name = "Raman Beta" ;
        rlprof_beta:units = "1/(m sr)" ;
        rlprof_beta:dpl_py_binding = "rlprofaerosol.beta" ;
    float rlprof_beta_error(time, altitude) ;
        rlprof_beta_error:long_name = "Uncertainty in calibrated aerosol volume backscatter coefficient" ;
        rlprof_beta_error:units = "1/(m sr)" ;
        rlprof_beta_error:dpl_py_binding = "rlprofaerosol.beta_error" ;
    float rlprof_ext_n2(time, altitude) ;
        rlprof_ext_n2:long_name = "Raman Aerosol N2 Extinction" ;
        rlprof_ext_n2:units = "1/m" ;
        rlprof_ext_n2:dpl_py_binding = "rlprofaerosol.extinction_n2" ;
    float rlprof_ext_n2_error(time, altitude) ;
        rlprof_ext_n2_error:long_name = "Uncertainty in aerosol extinction from N2" ;
        rlprof_ext_n2_error:units = "1/m" ;
        rlprof_ext_n2_error:dpl_py_binding = "rlprofaerosol.beta_error" ;
    float rlprof_bscat(time, altitude) ;
        rlprof_bscat:long_name = "Raman Aerosol Backscatter Extinction" ;
        rlprof_bscat:units = "1/m" ;
        rlprof_bscat:dpl_py_binding = "rlprofaerosol.extinction_bscat" ;
    float rlprof_bscat_error(time, altitude) ;
        rlprof_bscat_error:long_name = "Uncertainty in aerosol extinction from backscatter" ;
        rlprof_bscat_error:units = "1/m" ;
        rlprof_bscat_error:dpl_py_binding = "rlprofaerosol.extinction_bscat_error" ;
    float rlprof_sa(time, altitude) ;
        rlprof_sa:long_name = "Raman Extinction to Backscatter Ratio" ;
        rlprof_sa:units = "sr" ;
        rlprof_sa:dpl_py_binding = "rlprofaerosol.extinction_to_backscatter_ratio" ;
    float rlprof_sa_error(time, altitude) ;
        rlprof_sa_error:long_name = "Uncertainty in extinction to backscatter ratio" ;
        rlprof_sa_error:units = "sr" ;
        rlprof_sa_error:dpl_py_binding = "rlprofaerosol.extinction_to_backscatter_ratio_error" ;
    float rlprof_dep(time, altitude) ;
        rlprof_dep:long_name = "Raman Linear Depolarization" ;
        rlprof_dep:units = "percent" ;
        rlprof_dep:dpl_py_binding = "rlprofaerosol.linear_depol" ;
    float rlprof_dep_error(time, altitude) ;
        rlprof_dep_error:long_name = "Uncertainty in linear depolarization ratio" ;
        rlprof_dep_error:units = "unitless" ;
        rlprof_dep_error:dpl_py_binding = "rlprofaerosol.linear_depol_error" ;
        
    float rlprof_asr_profile(profile_time, altitude) ;
        rlprof_asr_profile:long_name = "Raman Aerosol Scattering Ratio" ;
        rlprof_asr_profile:units = "unitless" ;
        rlprof_asr_profile:dpl_py_binding = "rlprofaerosol_profile.aerosol_backscatter_ratio" ;
    float rlprof_asr_error_profile(profile_time, altitude) ;
        rlprof_asr_error_profile:long_name = "Uncertainty in calibrated aerosol scattering ratio" ;
        rlprof_asr_error_profile:units = "unitless" ;
        rlprof_asr_error_profile:dpl_py_binding = "rlprofaerosol_profile.aerosol_backscatter_ratio_error" ;
    float rlprof_beta_profile(profile_time, altitude) ;
        rlprof_beta_profile:long_name = "Raman Beta" ;
        rlprof_beta_profile:units = "1/(m sr)" ;
        rlprof_beta_profile:dpl_py_binding = "rlprofaerosol_profile.beta" ;
    float rlprof_beta_error_profile(profile_time, altitude) ;
        rlprof_beta_error_profile:long_name = "Uncertainty in calibrated aerosol volume backscatter coefficient" ;
        rlprof_beta_error_profile:units = "1/(m sr)" ;
        rlprof_beta_error_profile:dpl_py_binding = "rlprofaerosol_profile.beta_error" ;
    float rlprof_ext_n2_profile(profile_time, altitude) ;
        rlprof_ext_n2_profile:long_name = "Raman Aerosol N2 Extinction" ;
        rlprof_ext_n2_profile:units = "1/m" ;
        rlprof_ext_n2_profile:dpl_py_binding = "rlprofaerosol_profile.extinction_n2" ;
    float rlprof_ext_n2_error_profile(profile_time, altitude) ;
        rlprof_ext_n2_error_profile:long_name = "Uncertainty in aerosol extinction from N2" ;
        rlprof_ext_n2_error_profile:units = "1/m" ;
        rlprof_ext_n2_error_profile:dpl_py_binding = "rlprofaerosol_profile.beta_error" ;
    float rlprof_bscat_profile(profile_time, altitude) ;
        rlprof_bscat_profile:long_name = "Raman Aerosol Backscatter Extinction" ;
        rlprof_bscat_profile:units = "1/m" ;
        rlprof_bscat_profile:dpl_py_binding = "rlprofaerosol_profile.extinction_bscat" ;
    float rlprof_bscat_error_profile(profile_time, altitude) ;
        rlprof_bscat_error_profile:long_name = "Uncertainty in aerosol extinction from backscatter" ;
        rlprof_bscat_error_profile:units = "1/m" ;
        rlprof_bscat_error_profile:dpl_py_binding = "rlprofaerosol_profile.extinction_bscat_error" ;
    float rlprof_sa_profile(profile_time, altitude) ;
        rlprof_sa_profile:long_name = "Raman Extinction to Backscatter Ratio" ;
        rlprof_sa_profile:units = "sr" ;
        rlprof_sa_profile:dpl_py_binding = "rlprofaerosol_profile.extinction_to_backscatter_ratio" ;
    float rlprof_sa_error_profile(profile_time, altitude) ;
        rlprof_sa_error_profile:long_name = "Uncertainty in extinction to backscatter ratio" ;
        rlprof_sa_error_profile:units = "sr" ;
        rlprof_sa_error_profile:dpl_py_binding = "rlprofaerosol_profile.extinction_to_backscatter_ratio_error" ;
    float rlprof_dep_profile(profile_time, altitude) ;
        rlprof_dep_profile:long_name = "Raman Linear Depolarization" ;
        rlprof_dep_profile:units = "percent" ;
        rlprof_dep_profile:dpl_py_binding = "rlprofaerosol_profile.linear_depol" ;
    float rlprof_dep_error_profile(profile_time, altitude) ;
        rlprof_dep_error_profile:long_name = "Uncertainty in linear depolarization ratio" ;
        rlprof_dep_error_profile:units = "unitless" ;
        rlprof_dep_error_profile:dpl_py_binding = "rlprofaerosol_profile.linear_depol_error" ;

    float uw_rl_asr(time, altitude) ;
        uw_rl_asr:long_name = "UW-Computed Raman Aerosol Scattering Ratio" ;
        uw_rl_asr:units = "unitless" ;
        uw_rl_asr:dpl_py_binding = "raman_inv.aerosol_backscatter_ratio" ;
    float uw_rl_beta_r_355(altitude) ;
        uw_rl_beta_r_355:long_name = "UW-Computed Raman Beta 355nm" ;
        uw_rl_beta_r_355:units = "1/(m sr)" ;
        uw_rl_beta_r_355:dpl_py_binding = "raman_inv.beta_r_355" ;
    float uw_rl_beta_r_387(altitude) ;
        uw_rl_beta_r_387:long_name = "UW-Computed Raman Beta 387nm" ;
        uw_rl_beta_r_387:units = "1/(m sr)" ;
        uw_rl_beta_r_387:dpl_py_binding = "raman_inv.beta_r_387" ;
    float uw_rl_ext(time, altitude) ;
        uw_rl_ext:long_name = "UW-Computed Raman Extinction" ;
        uw_rl_ext:units = "" ;
        uw_rl_ext:dpl_py_binding = "raman_inv.extinction" ;
    float uw_rl_extaer(time, altitude) ;
        uw_rl_extaer:long_name = "UW-Computed Raman Aerosol Extinction" ;
        uw_rl_extaer:units = "" ;
        uw_rl_extaer:dpl_py_binding = "raman_inv.extinction_aerosol" ;
    float uw_rl_bscat(time, altitude) ;
        uw_rl_bscat:long_name = "UW-Computed Raman Aerosol Backscatter" ;
        uw_rl_bscat:units = "" ;
        uw_rl_bscat:dpl_py_binding = "raman_inv.beta_a_backscat" ;
    float uw_rl_intbscat(time, altitude) ;
        uw_rl_intbscat:long_name = "UW-Computed Raman Integrated Backscatter" ;
        uw_rl_intbscat:units = "" ;
        uw_rl_intbscat:dpl_py_binding = "raman_inv.integrated_backscatter" ;
    float uw_rl_dep(time, altitude) ;
        uw_rl_dep:long_name = "UW-Computed Raman Linear Depolarization" ;
        uw_rl_dep:units = "percent" ;
        uw_rl_dep:dpl_py_binding = "raman_inv.linear_depol" ;
    float uw_rl_od(time, altitude) ;
        uw_rl_od:long_name = "UW-Computed Raman Optical Depth" ;
        uw_rl_od:units = "" ;
        uw_rl_od:dpl_py_binding = "raman_inv.optical_depth" ;
    float uw_rl_p180(time, altitude) ;
        uw_rl_p180:long_name = "UW-Computed Raman P180" ;
        uw_rl_p180:units = "" ;
        uw_rl_p180:dpl_py_binding = "raman_inv.p180" ;

    float uw_rl_asr_profile(profile_time, altitude) ;
        uw_rl_asr_profile:long_name = "UW-Computed Raman Aerosol Scattering Ratio" ;
        uw_rl_asr_profile:units = "unitless" ;
        uw_rl_asr_profile:dpl_py_binding = "raman_profile.inv.aerosol_backscatter_ratio" ;
    float uw_rl_ext_profile(profile_time, altitude) ;
        uw_rl_ext_profile:long_name = "UW-Computed Raman Extinction" ;
        uw_rl_ext_profile:units = "" ;
        uw_rl_ext_profile:dpl_py_binding = "raman_profile.inv.extinction" ;
    float uw_rl_extaer_profile(profile_time, altitude) ;
        uw_rl_extaer_profile:long_name = "UW-Computed Raman Aerosol Extinction" ;
        uw_rl_extaer_profile:units = "" ;
        uw_rl_extaer_profile:dpl_py_binding = "raman_profile.inv.extinction_aerosol" ;
    float uw_rl_bscat_profile(profile_time, altitude) ;
        uw_rl_bscat_profile:long_name = "UW-Computed Raman Aerosol Backscatter" ;
        uw_rl_bscat_profile:units = "" ;
        uw_rl_bscat_profile:dpl_py_binding = "raman_profile.inv.beta_a_backscat" ;
    float uw_rl_intbscat_profile(profile_time, altitude) ;
        uw_rl_intbscat_profile:long_name = "UW-Computed Raman Integrated Backscatter" ;
        uw_rl_intbscat_profile:units = "" ;
        uw_rl_intbscat_profile:dpl_py_binding = "raman_profile.inv.integrated_backscatter" ;
    float uw_rl_dep_profile(profile_time, altitude) ;
        uw_rl_dep_profile:long_name = "UW-Computed Raman Linear Depolarization" ;
        uw_rl_dep_profile:units = "percent" ;
        uw_rl_dep_profile:dpl_py_binding = "raman_profile.inv.linear_depol" ;
    float uw_rl_od_profile(profile_time, altitude) ;
        uw_rl_od_profile:long_name = "UW-Computed Raman Optical Depth" ;
        uw_rl_od_profile:units = "" ;
        uw_rl_od_profile:dpl_py_binding = "raman_profile.inv.optical_depth" ;
    float uw_rl_p180_profile(profile_time, altitude) ;
        uw_rl_p180_profile:long_name = "UW-Computed Raman P180" ;
        uw_rl_p180_profile:units = "" ;
        uw_rl_p180_profile:dpl_py_binding = "raman_profile.inv.p180" ;

        float scattering_ratio_e_n2(time, altitude) ;
                scattering_ratio_e_n2:long_name = "Scattering ratio derived from the high elastic and nitrogen channels" ;
                scattering_ratio_e_n2:units = "unitless" ;
                scattering_ratio_e_n2:dpl_py_binding = "rlproffex1thor.scattering_ratio_e_n2" ;
        float scattering_ratio_e_n2_uncertainty(time, altitude, uncertainty) ;
                scattering_ratio_e_n2_uncertainty:long_name = "Uncertainty in scattering_ratio_e_n2" ;
                scattering_ratio_e_n2_uncertainty:units = "unitless" ;
                scattering_ratio_e_n2_uncertainty:comment = "Random: signal noise, calibration. Maximum systematic: weight, overlap, calibration" ;
                scattering_ratio_e_n2_uncertainty:dpl_py_binding = "rlproffex1thor.scattering_ratio_e_n2_uncertainty" ;
        float depolarization_ratio(time, altitude) ;
                depolarization_ratio:long_name = "Volume linear depolarization ratio" ;
                depolarization_ratio:units = "%" ;
                depolarization_ratio:comment = "Beam perpendicular component divided by the beam parallel component" ;
                depolarization_ratio:dpl_py_binding = "rlproffex1thor.depolarization_ratio" ;
        float depolarization_ratio_uncertainty(time, altitude, uncertainty) ;
                depolarization_ratio_uncertainty:long_name = "Uncertainty in depolarization_ratio" ;
                depolarization_ratio_uncertainty:units = "unitless" ;
                depolarization_ratio_uncertainty:comment = "Random: signal noise, misalignment angle. Maximum systematic: weight, misalignment angle" ;
                depolarization_ratio_uncertainty:dpl_py_binding = "rlproffex1thor.depolarization_ratio_uncertainty" ;
        float scattering_ratio_e(time, altitude) ;
                scattering_ratio_e:long_name = "Scattering ratio derived from the high elastic channels" ;
                scattering_ratio_e:units = "unitless" ;
                scattering_ratio_e:dpl_py_binding = "rlproffex1thor.scattering_ratio_e" ;
        double scattering_ratio_e_uncertainty(time, altitude, uncertainty) ;
                scattering_ratio_e_uncertainty:long_name = "Uncertainty in scattering_ratio_e" ;
                scattering_ratio_e_uncertainty:units = "unitless" ;
                scattering_ratio_e_uncertainty:comment = "Random: signal noise, calibration. Maximum systematic: weight, overlap, calibration" ;
                scattering_ratio_e_uncertainty:dpl_py_binding = "rlproffex1thor.scattering_ratio_e_uncertainty" ;
        float scattering_ratio_e_n2_low(time, altitude) ;
                scattering_ratio_e_n2_low:long_name = "Scattering ratio derived from the low elastic and nitrogen channels" ;
                scattering_ratio_e_n2_low:units = "unitless" ;
                scattering_ratio_e_n2_low:dpl_py_binding = "rlproffex1thor.scattering_ratio_e_n2_low" ;
        float scattering_ratio_e_n2_low_uncertainty(time, altitude, uncertainty) ;
                scattering_ratio_e_n2_low_uncertainty:long_name = "Uncertainty in scattering_ratio_e_n2_low" ;
                scattering_ratio_e_n2_low_uncertainty:units = "unitless" ;
                scattering_ratio_e_n2_low_uncertainty:comment = "Random: signal noise, calibration. Maximum systematic: calibration" ;
                scattering_ratio_e_n2_low_uncertainty:dpl_py_binding = "rlproffex1thor.scattering_ratio_e_n2_low_uncertainty" ;
        float particulate_backscatter_be(time, altitude) ;
                particulate_backscatter_be:long_name = "Best-estimate of the particulate backscatter coefficient" ;
                particulate_backscatter_be:units = "1/(m sr)" ;
                particulate_backscatter_be:comment = "Combination of: scattering_ratio_e_n2 + scattering_ratio_e_n2_low + Bp_el_beS as noted in extinction_flag" ;
                particulate_backscatter_be:dpl_py_binding = "rlproffex1thor.particulate_backscatter_be" ;
        float particulate_backscatter_be_uncertainty(time, altitude, uncertainty) ;
                particulate_backscatter_be_uncertainty:long_name = "Uncertainty in particulate_backscatter_be" ;
                particulate_backscatter_be_uncertainty:units = "1/(m sr)" ;
                particulate_backscatter_be_uncertainty:comment = "Random: scattering_ratio_e_n2_uncertainty scattering_ratio_e_n2_low_uncertainty Bp_el_beS_uncertainty. Maximum systematic: scattering_ratio_e_n2_uncertainty scattering_ratio_e_n2_low_uncertainty Bp_el_beS_uncertainty" ;
                particulate_backscatter_be_uncertainty:dpl_py_binding = "rlproffex1thor.particulate_backscatter_be_uncertainty" ;
        float lidar_ratio_be(time, altitude) ;
                lidar_ratio_be:long_name = "Best-estimate of the lidar ratio" ;
                lidar_ratio_be:units = "sr" ;
                lidar_ratio_be:comment = "Combination of: lidar_ratio_e_n2_low + lidar_ratio_e_n2 + interpolated + transmission-loss + profile/object/daily averaged + assumed lidar ratios as noted in extinction_flag" ;
                lidar_ratio_be:dpl_py_binding = "rlproffex1thor.lidar_ratio_be" ;
        float lidar_ratio_be_uncertainty(time, altitude, uncertainty) ;
                lidar_ratio_be_uncertainty:long_name = "Uncertainty in lidar_ratio_be" ;
                lidar_ratio_be_uncertainty:units = "sr" ;
                lidar_ratio_be_uncertainty:comment = "Random: signal noise, calibration, averaged lidar ratio. Maximum systematic: overlap, calibration, assumed lidar ratio, transmission optical depth, averaged lidar ratio" ;
                lidar_ratio_be_uncertainty:dpl_py_binding = "rlproffex1thor.lidar_ratio_be_uncertainty" ;
        float extinction_be(time, altitude) ;
                extinction_be:long_name = "Best-estimate of the particulate extinction coefficient" ;
                extinction_be:units = "1/m" ;
                extinction_be:comment = "particulate_backscatter_be * lidar_ratio_be" ;
                extinction_be:dpl_py_binding = "rlproffex1thor.extinction_be" ;
        float extinction_be_uncertainty(time, altitude, uncertainty) ;
                extinction_be_uncertainty:long_name = "Uncertainty in extinction_be" ;
                extinction_be_uncertainty:units = "1/m" ;
                extinction_be_uncertainty:comment = "Random: particulate_backscatter_be lidar_ratio_be. Maximum systematic: particulate_backscatter_be lidar_ratio_be" ;
                extinction_be_uncertainty:dpl_py_binding = "rlproffex1thor.extinction_be_uncertainty" ;
        float lidar_ratio_be_no_smooth(time, altitude) ;
                lidar_ratio_be_no_smooth:long_name = "Best-estimate of the lidar ratio without smoothing the transitions between sources" ;
                lidar_ratio_be_no_smooth:units = "sr" ;
                lidar_ratio_be_no_smooth:dpl_py_binding = "rlproffex1thor.lidar_ratio_be_no_smooth" ;
        float particulate_backscatter_be_no_smooth(time, altitude) ;
                particulate_backscatter_be_no_smooth:long_name = "Best-estimate particulate backscatter coefficient without smoothing the transitions between sources" ;
                particulate_backscatter_be_no_smooth:units = "1/(m sr)" ;
                particulate_backscatter_be_no_smooth:dpl_py_binding = "rlproffex1thor.particulate_backscatter_be_no_smooth" ;
        float particulate_backscatter_e_n2(time, altitude) ;
                particulate_backscatter_e_n2:long_name = "Particulate backscatter coefficient calculated from scattering_ratio_e_n2" ;
                particulate_backscatter_e_n2:units = "1/(m sr)" ;
                particulate_backscatter_e_n2:dpl_py_binding = "rlproffex1thor.particulate_backscatter_e_n2" ;
        float particulate_backscatter_n2_uncertainty(time, altitude, uncertainty) ;
                particulate_backscatter_n2_uncertainty:long_name = "Uncertainty in particulate_backscatter_e_n2" ;
                particulate_backscatter_n2_uncertainty:units = "1/(m sr)" ;
                particulate_backscatter_n2_uncertainty:comment = "Random: scattering_ratio_e_n2_uncertainty. Maximum systematic: scattering_ratio_e_n2_uncertainty" ;
                particulate_backscatter_n2_uncertainty:dpl_py_binding = "rlproffex1thor.particulate_backscatter_n2_uncertainty" ;
        float particulate_backscatter_e_n2_low(time, altitude) ;
                particulate_backscatter_e_n2_low:long_name = "Particulate backscatter coefficient calculated from scattering_ratio_e_n2_low" ;
                particulate_backscatter_e_n2_low:units = "1/(m sr)" ;
                particulate_backscatter_e_n2_low:dpl_py_binding = "rlproffex1thor.particulate_backscatter_e_n2_low" ;
        float particulate_backscatter_n2_low_uncertainty(time, altitude, uncertainty) ;
                particulate_backscatter_n2_low_uncertainty:long_name = "Uncertainty in particulate_backscatter_n2_low" ;
                particulate_backscatter_n2_low_uncertainty:units = "1/(m sr)" ;
                particulate_backscatter_n2_low_uncertainty:comment = "Random: scattering_ratio_e_n2_low_uncertainty. Maximum systematic: scattering_ratio_e_n2_low_uncertainty" ;
                particulate_backscatter_n2_low_uncertainty:dpl_py_binding = "rlproffex1thor.particulate_backscatter_n2_low_uncertainty" ;
        float particulate_backscatter_e_beS(time, altitude) ;
                particulate_backscatter_e_beS:long_name = "Particulate backscatter coefficient from the high elastic channels using the best-estimate lidar ratios" ;
                particulate_backscatter_e_beS:units = "1/(m sr)" ;
                particulate_backscatter_e_beS:comment = "Fernald solution using lidar_ratio_be" ;
                particulate_backscatter_e_beS:dpl_py_binding = "rlproffex1thor.particulate_backscatter_e_beS" ;
        float particulate_backscatter_e_beS_uncertainty(time, altitude, uncertainty) ;
                particulate_backscatter_e_beS_uncertainty:long_name = "Uncertainty in particulate_backscatter_e_beS" ;
                particulate_backscatter_e_beS_uncertainty:units = "1/(m sr)" ;
                particulate_backscatter_e_beS_uncertainty:comment = "Random: signal noise, lidar_ratio_be_uncertainty. Maximum systematic: lidar_ratio_be_uncertainty" ;
                particulate_backscatter_e_beS_uncertainty:dpl_py_binding = "rlproffex1thor.particulate_backscatter_e_beS_uncertainty" ;
        float particulate_backscatter_e(time, altitude) ;
                particulate_backscatter_e:long_name = "Particulate backscatter coefficient from the high elastic channels" ;
                particulate_backscatter_e:units = "1/(m sr)" ;
                particulate_backscatter_e:comment = "Fernald solution using the lidar ratios given in lidar_ratio_e" ;
                particulate_backscatter_e:dpl_py_binding = "rlproffex1thor.particulate_backscatter_e" ;
        float particulate_backscatter_e_uncertainty(time, altitude, uncertainty) ;
                particulate_backscatter_e_uncertainty:long_name = "Uncertainty in particulate_backscatter_e" ;
                particulate_backscatter_e_uncertainty:units = "1/(m sr)" ;
                particulate_backscatter_e_uncertainty:comment = "Random: signal noise. Maximum systematic: assumed lidar ratio, transmission optical depth" ;
                particulate_backscatter_e_uncertainty:dpl_py_binding = "rlproffex1thor.particulate_backscatter_e_uncertainty" ;
        float lidar_ratio_e_n2(time, altitude) ;
                lidar_ratio_e_n2:long_name = "Lidar ratio from the high nitrogen channel extinction and particulate_backscatter_e_n2" ;
                lidar_ratio_e_n2:units = "sr" ;
                lidar_ratio_e_n2:comment = "Determined at various amounts of smoothing as noted in extinction_flag" ;
                lidar_ratio_e_n2:dpl_py_binding = "rlproffex1thor.lidar_ratio_e_n2" ;
        float lidar_ratio_e_n2_uncertainty(time, altitude, uncertainty) ;
                lidar_ratio_e_n2_uncertainty:long_name = "Uncertainty lidar_ratio_e_n2" ;
                lidar_ratio_e_n2_uncertainty:units = "sr" ;
                lidar_ratio_e_n2_uncertainty:comment = "Random: signal noise. Maximum systematic: N/A" ;
                lidar_ratio_e_n2_uncertainty:dpl_py_binding = "rlproffex1thor.lidar_ratio_e_n2_uncertainty" ;
        float lidar_ratio_e_n2_low(time, altitude) ;
                lidar_ratio_e_n2_low:long_name = "Lidar ratio from the low nitrogen channel extinction and particulate_backscatter_e_n2_low" ;
                lidar_ratio_e_n2_low:units = "sr" ;
                lidar_ratio_e_n2_low:comment = "Determined at various amounts of smoothing as noted in extinction_flag" ;
                lidar_ratio_e_n2_low:dpl_py_binding = "rlproffex1thor.lidar_ratio_e_n2_low" ;
        float lidar_ratio_e_n2_low_uncertainty(time, altitude, uncertainty) ;
                lidar_ratio_e_n2_low_uncertainty:long_name = "Uncertainty in lidar_ratio_e_n2_low" ;
                lidar_ratio_e_n2_low_uncertainty:units = "sr" ;
                lidar_ratio_e_n2_low_uncertainty:comment = "Random: signal noise. Maximum systematic: N/A" ;
                lidar_ratio_e_n2_low_uncertainty:dpl_py_binding = "rlproffex1thor.lidar_ratio_e_n2_low_uncertainty" ;
        float lidar_ratio_e(time, altitude) ;
                lidar_ratio_e:long_name = "Lidar ratio from the high elastic channels" ;
                lidar_ratio_e:units = "sr" ;
                lidar_ratio_e:comment = "Combination of assumed values based on feature type and values determined from the transmission-loss method" ;
                lidar_ratio_e:dpl_py_binding = "rlproffex1thor.lidar_ratio_e" ;
        float lidar_ratio_e_uncertainty(time, altitude, uncertainty) ;
                lidar_ratio_e_uncertainty:long_name = "Uncertainty in lidar_ratio_e" ;
                lidar_ratio_e_uncertainty:units = "sr" ;
                lidar_ratio_e_uncertainty:comment = "Random: signal noise. Maximum systematic: assumed lidar ratio, transmission optical depth" ;
                lidar_ratio_e_uncertainty:dpl_py_binding = "rlproffex1thor.lidar_ratio_e_uncertainty" ;
        float particulate_backscatter_be_noMS(time, altitude) ;
                particulate_backscatter_be_noMS:long_name = "Best-estimate of the particulate backscatter coefficient without accounting for multiple scattering effects" ;
                particulate_backscatter_be_noMS:units = "1/(m sr)" ;
                particulate_backscatter_be_noMS:comment = "Combination of: scattering_ratio_e_n2 + scattering_ratio_e_n2_low + Bp_el_beS as noted in extinction_flag" ;
                particulate_backscatter_be_noMS:dpl_py_binding = "rlproffex1thor.particulate_backscatter_be_noMS" ;
        float lidar_ratio_be_noMS(time, altitude) ;
                lidar_ratio_be_noMS:long_name = "Best-estimate of the lidar ratio without accounting for multiple scattering effects" ;
                lidar_ratio_be_noMS:units = "sr" ;
                lidar_ratio_be_noMS:comment = "Combination of: lidar_ratio_e_n2_low + lidar_ratio_e_n2 + interpolated + transmission-loss + profile/object/daily averaged + assumed lidar ratios as noted in extinction_flag" ;
                lidar_ratio_be_noMS:dpl_py_binding = "rlproffex1thor.lidar_ratio_be_noMS" ;
        float lidar_ratio_e_n2_noMS(time, altitude) ;
                lidar_ratio_e_n2_noMS:long_name = "Lidar ratio from the high nitrogen channel extinction and particulate_backscatter_e_n2 without accounting for multiple scattering effects" ;
                lidar_ratio_e_n2_noMS:units = "sr" ;
                lidar_ratio_e_n2_noMS:comment = "Determined at various amounts of smoothing as noted in extinction_flag" ;
                lidar_ratio_e_n2_noMS:dpl_py_binding = "rlproffex1thor.lidar_ratio_e_n2_noMS" ;
        float lidar_ratio_e_n2_low_noMS(time, altitude) ;
                lidar_ratio_e_n2_low_noMS:long_name = "Lidar ratio from the low nitrogen channel extinction and particulate_backscatter_e_n2_low without accounting for multiple scattering effects" ;
                lidar_ratio_e_n2_low_noMS:units = "sr" ;
                lidar_ratio_e_n2_low_noMS:comment = "Determined at various amounts of smoothing as noted in extinction_flag" ;
                lidar_ratio_e_n2_low_noMS:dpl_py_binding = "rlproffex1thor.lidar_ratio_e_n2_low_noMS" ;
        float lidar_ratio_e_noMS(time, altitude) ;
                lidar_ratio_e_noMS:long_name = "Lidar ratio from the high elastic channels without accounting for multiple scattering effects" ;
                lidar_ratio_e_noMS:units = "sr" ;
                lidar_ratio_e_noMS:comment = "Combination of assumed values based on feature type and values determined from the transmission-loss method" ;
                lidar_ratio_e_noMS:dpl_py_binding = "rlproffex1thor.lidar_ratio_e_noMS" ;

        float scattering_ratio_e_n2_profile(profile_time, altitude) ;
                scattering_ratio_e_n2_profile:long_name = "Scattering ratio derived from the high elastic and nitrogen channels" ;
                scattering_ratio_e_n2_profile:units = "unitless" ;
                scattering_ratio_e_n2_profile:dpl_py_binding = "rlproffex1thor_profile.scattering_ratio_e_n2" ;
        float scattering_ratio_e_n2_uncertainty_profile(profile_time, altitude, uncertainty) ;
                scattering_ratio_e_n2_uncertainty_profile:long_name = "Uncertainty in scattering_ratio_e_n2" ;
                scattering_ratio_e_n2_uncertainty_profile:units = "unitless" ;
                scattering_ratio_e_n2_uncertainty_profile:comment = "Random: signal noise, calibration. Maximum systematic: weight, overlap, calibration" ;
                scattering_ratio_e_n2_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.scattering_ratio_e_n2_uncertainty" ;
        float depolarization_ratio_profile(profile_time, altitude) ;
                depolarization_ratio_profile:long_name = "Volume linear depolarization ratio" ;
                depolarization_ratio_profile:units = "%" ;
                depolarization_ratio_profile:comment = "Beam perpendicular component divided by the beam parallel component" ;
                depolarization_ratio_profile:dpl_py_binding = "rlproffex1thor_profile.depolarization_ratio" ;
        float depolarization_ratio_uncertainty_profile(profile_time, altitude, uncertainty) ;
                depolarization_ratio_uncertainty_profile:long_name = "Uncertainty in depolarization_ratio" ;
                depolarization_ratio_uncertainty_profile:units = "unitless" ;
                depolarization_ratio_uncertainty_profile:comment = "Random: signal noise, misalignment angle. Maximum systematic: weight, misalignment angle" ;
                depolarization_ratio_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.depolarization_ratio_uncertainty" ;
        float scattering_ratio_e_profile(profile_time, altitude) ;
                scattering_ratio_e_profile:long_name = "Scattering ratio derived from the high elastic channels" ;
                scattering_ratio_e_profile:units = "unitless" ;
                scattering_ratio_e_profile:dpl_py_binding = "rlproffex1thor_profile.scattering_ratio_e" ;
        double scattering_ratio_e_uncertainty_profile(profile_time, altitude, uncertainty) ;
                scattering_ratio_e_uncertainty_profile:long_name = "Uncertainty in scattering_ratio_e" ;
                scattering_ratio_e_uncertainty_profile:units = "unitless" ;
                scattering_ratio_e_uncertainty_profile:comment = "Random: signal noise, calibration. Maximum systematic: weight, overlap, calibration" ;
                scattering_ratio_e_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.scattering_ratio_e_uncertainty" ;
        float scattering_ratio_e_n2_low_profile(profile_time, altitude) ;
                scattering_ratio_e_n2_low_profile:long_name = "Scattering ratio derived from the low elastic and nitrogen channels" ;
                scattering_ratio_e_n2_low_profile:units = "unitless" ;
                scattering_ratio_e_n2_low_profile:dpl_py_binding = "rlproffex1thor_profile.scattering_ratio_e_n2_low" ;
        float scattering_ratio_e_n2_low_uncertainty_profile(profile_time, altitude, uncertainty) ;
                scattering_ratio_e_n2_low_uncertainty_profile:long_name = "Uncertainty in scattering_ratio_e_n2_low" ;
                scattering_ratio_e_n2_low_uncertainty_profile:units = "unitless" ;
                scattering_ratio_e_n2_low_uncertainty_profile:comment = "Random: signal noise, calibration. Maximum systematic: calibration" ;
                scattering_ratio_e_n2_low_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.scattering_ratio_e_n2_low_uncertainty" ;
        float particulate_backscatter_be_profile(profile_time, altitude) ;
                particulate_backscatter_be_profile:long_name = "Best-estimate of the particulate backscatter coefficient" ;
                particulate_backscatter_be_profile:units = "1/(m sr)" ;
                particulate_backscatter_be_profile:comment = "Combination of: scattering_ratio_e_n2 + scattering_ratio_e_n2_low + Bp_el_beS as noted in extinction_flag" ;
                particulate_backscatter_be_profile:dpl_py_binding = "rlproffex1thor_profile.particulate_backscatter_be" ;
        float particulate_backscatter_be_uncertainty_profile(profile_time, altitude, uncertainty) ;
                particulate_backscatter_be_uncertainty_profile:long_name = "Uncertainty in particulate_backscatter_be" ;
                particulate_backscatter_be_uncertainty_profile:units = "1/(m sr)" ;
                particulate_backscatter_be_uncertainty_profile:comment = "Random: scattering_ratio_e_n2_uncertainty scattering_ratio_e_n2_low_uncertainty Bp_el_beS_uncertainty. Maximum systematic: scattering_ratio_e_n2_uncertainty scattering_ratio_e_n2_low_uncertainty Bp_el_beS_uncertainty" ;
                particulate_backscatter_be_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.particulate_backscatter_be_uncertainty" ;
        float lidar_ratio_be_profile(profile_time, altitude) ;
                lidar_ratio_be_profile:long_name = "Best-estimate of the lidar ratio" ;
                lidar_ratio_be_profile:units = "sr" ;
                lidar_ratio_be_profile:comment = "Combination of: lidar_ratio_e_n2_low + lidar_ratio_e_n2 + interpolated + transmission-loss + profile/object/daily averaged + assumed lidar ratios as noted in extinction_flag" ;
                lidar_ratio_be_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_be" ;
        float lidar_ratio_be_uncertainty_profile(profile_time, altitude, uncertainty) ;
                lidar_ratio_be_uncertainty_profile:long_name = "Uncertainty in lidar_ratio_be" ;
                lidar_ratio_be_uncertainty_profile:units = "sr" ;
                lidar_ratio_be_uncertainty_profile:comment = "Random: signal noise, calibration, averaged lidar ratio. Maximum systematic: overlap, calibration, assumed lidar ratio, transmission optical depth, averaged lidar ratio" ;
                lidar_ratio_be_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_be_uncertainty" ;
        float extinction_be_profile(profile_time, altitude) ;
                extinction_be_profile:long_name = "Best-estimate of the particulate extinction coefficient" ;
                extinction_be_profile:units = "1/m" ;
                extinction_be_profile:comment = "particulate_backscatter_be * lidar_ratio_be" ;
                extinction_be_profile:dpl_py_binding = "rlproffex1thor_profile.extinction_be" ;
        float extinction_be_uncertainty_profile(profile_time, altitude, uncertainty) ;
                extinction_be_uncertainty_profile:long_name = "Uncertainty in extinction_be" ;
                extinction_be_uncertainty_profile:units = "1/m" ;
                extinction_be_uncertainty_profile:comment = "Random: particulate_backscatter_be lidar_ratio_be. Maximum systematic: particulate_backscatter_be lidar_ratio_be" ;
                extinction_be_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.extinction_be_uncertainty" ;
        float lidar_ratio_be_no_smooth_profile(time, altitude) ;
                lidar_ratio_be_no_smooth_profile:long_name = "Best-estimate of the lidar ratio without smoothing the transitions between sources" ;
                lidar_ratio_be_no_smooth_profile:units = "sr" ;
                lidar_ratio_be_no_smooth_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_be_no_smooth" ;
        float particulate_backscatter_be_no_smooth_profile(profile_time, altitude) ;
                particulate_backscatter_be_no_smooth_profile:long_name = "Best-estimate particulate backscatter coefficient without smoothing the transitions between sources" ;
                particulate_backscatter_be_no_smooth_profile:units = "1/(m sr)" ;
                particulate_backscatter_be_no_smooth_profile:dpl_py_binding = "rlproffex1thor_profile.particulate_backscatter_be_no_smooth" ;
        float particulate_backscatter_e_n2_profile(profile_time, altitude) ;
                particulate_backscatter_e_n2_profile:long_name = "Particulate backscatter coefficient calculated from scattering_ratio_e_n2" ;
                particulate_backscatter_e_n2_profile:units = "1/(m sr)" ;
                particulate_backscatter_e_n2_profile:dpl_py_binding = "rlproffex1thor_profile.particulate_backscatter_e_n2" ;
        float particulate_backscatter_n2_uncertainty_profile(profile_time, altitude, uncertainty) ;
                particulate_backscatter_n2_uncertainty_profile:long_name = "Uncertainty in particulate_backscatter_e_n2" ;
                particulate_backscatter_n2_uncertainty_profile:units = "1/(m sr)" ;
                particulate_backscatter_n2_uncertainty_profile:comment = "Random: scattering_ratio_e_n2_uncertainty. Maximum systematic: scattering_ratio_e_n2_uncertainty" ;
                particulate_backscatter_n2_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.particulate_backscatter_n2_uncertainty" ;
        float particulate_backscatter_e_n2_low_profile(profile_time, altitude) ;
                particulate_backscatter_e_n2_low_profile:long_name = "Particulate backscatter coefficient calculated from scattering_ratio_e_n2_low" ;
                particulate_backscatter_e_n2_low_profile:units = "1/(m sr)" ;
                particulate_backscatter_e_n2_low_profile:dpl_py_binding = "rlproffex1thor_profile.particulate_backscatter_e_n2_low" ;
        float particulate_backscatter_n2_low_uncertainty_profile(profile_time, altitude, uncertainty) ;
                particulate_backscatter_n2_low_uncertainty_profile:long_name = "Uncertainty in particulate_backscatter_n2_low" ;
                particulate_backscatter_n2_low_uncertainty_profile:units = "1/(m sr)" ;
                particulate_backscatter_n2_low_uncertainty_profile:comment = "Random: scattering_ratio_e_n2_low_uncertainty. Maximum systematic: scattering_ratio_e_n2_low_uncertainty" ;
                particulate_backscatter_n2_low_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.particulate_backscatter_n2_low_uncertainty" ;
        float particulate_backscatter_e_beS_profile(profile_time, altitude) ;
                particulate_backscatter_e_beS_profile:long_name = "Particulate backscatter coefficient from the high elastic channels using the best-estimate lidar ratios" ;
                particulate_backscatter_e_beS_profile:units = "1/(m sr)" ;
                particulate_backscatter_e_beS_profile:comment = "Fernald solution using lidar_ratio_be" ;
                particulate_backscatter_e_beS_profile:dpl_py_binding = "rlproffex1thor_profile.particulate_backscatter_e_beS" ;
        float particulate_backscatter_e_beS_uncertainty_profile(profile_time, altitude, uncertainty) ;
                particulate_backscatter_e_beS_uncertainty_profile:long_name = "Uncertainty in particulate_backscatter_e_beS" ;
                particulate_backscatter_e_beS_uncertainty_profile:units = "1/(m sr)" ;
                particulate_backscatter_e_beS_uncertainty_profile:comment = "Random: signal noise, lidar_ratio_be_uncertainty. Maximum systematic: lidar_ratio_be_uncertainty" ;
                particulate_backscatter_e_beS_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.particulate_backscatter_e_beS_uncertainty" ;
        float particulate_backscatter_e_profile(profile_time, altitude) ;
                particulate_backscatter_e_profile:long_name = "Particulate backscatter coefficient from the high elastic channels" ;
                particulate_backscatter_e_profile:units = "1/(m sr)" ;
                particulate_backscatter_e_profile:comment = "Fernald solution using the lidar ratios given in lidar_ratio_e" ;
                particulate_backscatter_e_profile:dpl_py_binding = "rlproffex1thor_profile.particulate_backscatter_e" ;
        float particulate_backscatter_e_uncertainty_profile(profile_time, altitude, uncertainty) ;
                particulate_backscatter_e_uncertainty_profile:long_name = "Uncertainty in particulate_backscatter_e" ;
                particulate_backscatter_e_uncertainty_profile:units = "1/(m sr)" ;
                particulate_backscatter_e_uncertainty_profile:comment = "Random: signal noise. Maximum systematic: assumed lidar ratio, transmission optical depth" ;
                particulate_backscatter_e_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.particulate_backscatter_e_uncertainty" ;
        float lidar_ratio_e_n2_profile(profile_time, altitude) ;
                lidar_ratio_e_n2_profile:long_name = "Lidar ratio from the high nitrogen channel extinction and particulate_backscatter_e_n2" ;
                lidar_ratio_e_n2_profile:units = "sr" ;
                lidar_ratio_e_n2_profile:comment = "Determined at various amounts of smoothing as noted in extinction_flag" ;
                lidar_ratio_e_n2_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_e_n2" ;
        float lidar_ratio_e_n2_uncertainty_profile(profile_time, altitude, uncertainty) ;
                lidar_ratio_e_n2_uncertainty_profile:long_name = "Uncertainty lidar_ratio_e_n2" ;
                lidar_ratio_e_n2_uncertainty_profile:units = "sr" ;
                lidar_ratio_e_n2_uncertainty_profile:comment = "Random: signal noise. Maximum systematic: N/A" ;
                lidar_ratio_e_n2_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_e_n2_uncertainty" ;
        float lidar_ratio_e_n2_low_profile(profile_time, altitude) ;
                lidar_ratio_e_n2_low_profile:long_name = "Lidar ratio from the low nitrogen channel extinction and particulate_backscatter_e_n2_low" ;
                lidar_ratio_e_n2_low_profile:units = "sr" ;
                lidar_ratio_e_n2_low_profile:comment = "Determined at various amounts of smoothing as noted in extinction_flag" ;
                lidar_ratio_e_n2_low_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_e_n2_low" ;
        float lidar_ratio_e_n2_low_uncertainty_profile(profile_time, altitude, uncertainty) ;
                lidar_ratio_e_n2_low_uncertainty_profile:long_name = "Uncertainty in lidar_ratio_e_n2_low" ;
                lidar_ratio_e_n2_low_uncertainty_profile:units = "sr" ;
                lidar_ratio_e_n2_low_uncertainty_profile:comment = "Random: signal noise. Maximum systematic: N/A" ;
                lidar_ratio_e_n2_low_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_e_n2_low_uncertainty" ;
        float lidar_ratio_e_profile(profile_time, altitude) ;
                lidar_ratio_e_profile:long_name = "Lidar ratio from the high elastic channels" ;
                lidar_ratio_e_profile:units = "sr" ;
                lidar_ratio_e_profile:comment = "Combination of assumed values based on feature type and values determined from the transmission-loss method" ;
                lidar_ratio_e_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_e" ;
        float lidar_ratio_e_uncertainty_profile(profile_time, altitude, uncertainty) ;
                lidar_ratio_e_uncertainty_profile:long_name = "Uncertainty in lidar_ratio_e" ;
                lidar_ratio_e_uncertainty_profile:units = "sr" ;
                lidar_ratio_e_uncertainty_profile:comment = "Random: signal noise. Maximum systematic: assumed lidar ratio, transmission optical depth" ;
                lidar_ratio_e_uncertainty_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_e_uncertainty" ;
        float particulate_backscatter_be_noMS_profile(profile_time, altitude) ;
                particulate_backscatter_be_noMS_profile:long_name = "Best-estimate of the particulate backscatter coefficient without accounting for multiple scattering effects" ;
                particulate_backscatter_be_noMS_profile:units = "1/(m sr)" ;
                particulate_backscatter_be_noMS_profile:comment = "Combination of: scattering_ratio_e_n2 + scattering_ratio_e_n2_low + Bp_el_beS as noted in extinction_flag" ;
                particulate_backscatter_be_noMS_profile:dpl_py_binding = "rlproffex1thor_profile.particulate_backscatter_be_noMS" ;
        float lidar_ratio_be_noMS_profile(profile_time, altitude) ;
                lidar_ratio_be_noMS_profile:long_name = "Best-estimate of the lidar ratio without accounting for multiple scattering effects" ;
                lidar_ratio_be_noMS_profile:units = "sr" ;
                lidar_ratio_be_noMS_profile:comment = "Combination of: lidar_ratio_e_n2_low + lidar_ratio_e_n2 + interpolated + transmission-loss + profile/object/daily averaged + assumed lidar ratios as noted in extinction_flag" ;
                lidar_ratio_be_noMS_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_be_noMS" ;
        float lidar_ratio_e_n2_noMS_profile(profile_time, altitude) ;
                lidar_ratio_e_n2_noMS_profile:long_name = "Lidar ratio from the high nitrogen channel extinction and particulate_backscatter_e_n2 without accounting for multiple scattering effects" ;
                lidar_ratio_e_n2_noMS_profile:units = "sr" ;
                lidar_ratio_e_n2_noMS_profile:comment = "Determined at various amounts of smoothing as noted in extinction_flag" ;
                lidar_ratio_e_n2_noMS_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_e_n2_noMS" ;
        float lidar_ratio_e_n2_low_noMS_profile(profile_time, altitude) ;
                lidar_ratio_e_n2_low_noMS_profile:long_name = "Lidar ratio from the low nitrogen channel extinction and particulate_backscatter_e_n2_low without accounting for multiple scattering effects" ;
                lidar_ratio_e_n2_low_noMS_profile:units = "sr" ;
                lidar_ratio_e_n2_low_noMS_profile:comment = "Determined at various amounts of smoothing as noted in extinction_flag" ;
                lidar_ratio_e_n2_low_noMS_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_e_n2_low_noMS" ;
        float lidar_ratio_e_noMS_profile(profile_time, altitude) ;
                lidar_ratio_e_noMS_profile:long_name = "Lidar ratio from the high elastic channels without accounting for multiple scattering effects" ;
                lidar_ratio_e_noMS_profile:units = "sr" ;
                lidar_ratio_e_noMS_profile:comment = "Combination of assumed values based on feature type and values determined from the transmission-loss method" ;
                lidar_ratio_e_noMS_profile:dpl_py_binding = "rlproffex1thor_profile.lidar_ratio_e_noMS" ;

// global attributes:
        :dpl_py_template = "hsrl_nomenclature.cdl" ;
        :dpl_py_template_version = 20161111 ;
        :time_zone = "UTC" ;
}
