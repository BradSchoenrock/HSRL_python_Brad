netcdf out {
dimensions:
	time = UNLIMITED ;
	sweep = 1 ;
	range = 0 ;
	bin_range = 0;
	profile_time = 1;
	time_vector = 8 ;
	calibration = UNLIMITED ; 
	githash = 40;
	sondenamelength = 10 ;
	i2header = 1000 ;
	geoheader = 1000 ;
	apheader = 1000 ;
	aeri_btemp_wavenumber = 0 ;
	aeri_mean_rad_wavenumber_ch1 = 0 ;
	aeri_mean_rad_wavenumber_ch2 = 0 ;
	mwr_frequency = 0 ;
	string_length_short = 32;
variables:
	char time_coverage_start(string_length_short) ;
		time_coverage_start:standard_name = "data_volume_start_time_utc" ;
		time_coverage_start:comment = "ray times are relative to start time in secs" ;
	char time_coverage_end(string_length_short) ;
		time_coverage_end:standard_name = "data_volume_end_time_utc" ;
	short first_time(time_vector) ;
		first_time:long_name = "First Time in file" ;
		first_time:dpl_py_binding = "dne" ;
	double sonde_times(calibration) ;
		sonde_times:long_name = "Time of Temperature Profiles" ;
		sonde_times:description = "New raob data" ;
		sonde_times:dpl_py_binding = "sounding.times" ;
        sonde_times:dpl_py_type = "python_datetime" ;
	double sonde_longitude(calibration) ;
		sonde_longitude:long_name = "Longitude of Temperature Profiles" ;
		sonde_longitude:units = "degrees_east" ;
		sonde_longitude:description = "Sounding Longitude source" ;
		sonde_longitude:dpl_py_binding = "sounding.longitude" ;
	double sonde_latitude(calibration) ;
		sonde_latitude:long_name = "Latituide of Temperature Profiles" ;
		sonde_latitude:units = "degrees_north" ;
		sonde_latitude:description = "Sounding Latitude source" ;
		sonde_latitude:dpl_py_binding = "sounding.latitude" ;
	double new_cal_times(calibration) ;
		new_cal_times:long_name = "Time of Calibration Change" ;
		new_cal_times:description = "New raob or system calibration data triggered recalibration" ;
		new_cal_times:dpl_py_binding = "chunk_start_time" ;
        new_cal_times:dpl_py_type = "python_datetime" ;
	byte new_cal_trigger(calibration) ;
		new_cal_trigger:long_name = "Trigger of Calibration Change" ;
		new_cal_trigger:description = "reason for recalibration" ;
		new_cal_trigger:bit_0 = "radiosonde profile" ;
		new_cal_trigger:bit_1 = "i2 scan" ;
		new_cal_trigger:bit_2 = "geometry" ;
		new_cal_trigger:dpl_py_binding = "dne" ;
	short new_cal_offset(calibration) ;
		new_cal_offset:long_name = "Record Dimension equivalent Offset" ;
		new_cal_offset:min_value = 0 ;
		new_cal_offset:dpl_py_binding = "dne" ;
	float top_alt_sounding(calibration) ;
		top_alt_sounding:long_name = "Sounding Maximum Altitude" ;
		top_alt_sounding:units = "meters" ;
		top_alt_sounding:dpl_py_binding = "sounding.top" ;
	float temperature_profile(time, range) ;
		temperature_profile:long_name = "Raob Temperature Profile" ;
		temperature_profile:description = "Temperature interpolated to requested altitude resolution" ;
		temperature_profile:units = "degrees Kelvin" ;
		temperature_profile:dpl_py_binding = "rs_inv.temps" ;
	float pressure_profile(time, range) ;
		pressure_profile:long_name = "Raob pressure Profile" ;
		pressure_profile:description = "Pressure interpolated to requested altitude resolution" ;
		pressure_profile:units = "hectopascals" ;
		pressure_profile:dpl_py_binding = "rs_inv.pressures" ;
	float dewpoint_profile(time, range) ;
		dewpoint_profile:long_name = "Raob Dewpoint Temperature Profile" ;
		dewpoint_profile:description = "Dewpoint interpolated to requested altitude resolution" ;
		dewpoint_profile:units = "degrees Kelvin" ;
		dewpoint_profile:missing_value = 9.96920996838687e+36 ;
		dewpoint_profile:dpl_py_binding = "rs_inv.dew_points" ;
	float windspeed_profile(time, range) ;
		windspeed_profile:long_name = "Raob Wind Speed Profile" ;
		windspeed_profile:description = "Speeds interpolated to requested altitude resolution" ;
		windspeed_profile:units = "m/s" ;
		windspeed_profile:missing_value = 9.96920996838687e+36 ;
		windspeed_profile:dpl_py_binding = "rs_inv.wind_spd" ;
	float winddir_profile(time, range) ;
		winddir_profile:long_name = "Raob Wind Direction Profile" ;
		winddir_profile:description = "Directions interpolated to requested altitude resolution" ;
		winddir_profile:units = "degrees" ;
		winddir_profile:missing_value = 9.96920996838687e+36 ;
		winddir_profile:dpl_py_binding = "rs_inv.wind_dir" ;
	char calibration_version(calibration, githash) ;
		calibration_version:long_name = "Calibration Tables GIT Version" ;
		calibration_version:dpl_py_binding = "gitversion" ;
	char raob_station(calibration, sondenamelength) ;
		raob_station:long_name = "Radiosonde Station ID" ;
		raob_station:dpl_py_binding = "sounding.sounding_id" ;
	char i2_txt_header(calibration, i2header) ;
		i2_txt_header:long_name = "i2_scan_file_text_info" ;
		i2_txt_header:description = "Contains name of file used to compute calibration" ;
		i2_txt_header:dpl_py_binding = "rs_cal.i2scan.header" ;
	char geo_txt_header(calibration, geoheader) ;
		geo_txt_header:long_name = "geometric_correction_file_txt_header." ;
		geo_txt_header:dpl_py_binding = "rs_cal.geo.header" ;
	char ap_txt_header(calibration, apheader) ;
		ap_txt_header:long_name = "afterpulse_correction_file_txt_header." ;
		ap_txt_header:dpl_py_binding = "rs_cal.afterpulse.header" ;
	float Cmc(calibration, range) ;
		Cmc:long_name = "Molecular in Combined Calibration" ;
		Cmc:dpl_py_binding = "rs_Cxx.Cmc" ;
	float Cmm(calibration, range) ;
		Cmm:long_name = "Molecular in Molecular Calibration" ;
		Cmm:dpl_py_binding = "rs_Cxx.Cmm" ;
	float Cam(calibration) ;
		Cam:long_name = "Aerosol in Molecular Calibration" ;
		Cam:dpl_py_binding = "rs_Cxx.Cam" ;
	float Cmm_i2a(calibration, range) ;
		Cmm_i2a:long_name = "Molecular in Molecular Calibration" ;
		Cmm_i2a:dpl_py_binding = "rs_Cxx.Cmm_i2a" ;
	short last_time(time_vector) ;
		last_time:long_name = "Last Time in file" ;
		last_time:dpl_py_binding = "dne" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time in seconds since volume start" ;
		time:units = "seconds since 2006-10-23 18:19:59 UTC" ;
		time:comment = "times are relative to the volume start_time" ;
		time:dpl_py_binding = "rs_inv.times" ;
		time:dpl_py_type = "python_datetime" ;
	double mean_time(time) ;
		mean_time:long_name = "Mean Time" ;
		mean_time:units = "seconds since 2006-10-23 18:19:59 UTC" ;
		mean_time:dpl_py_binding = "rs_mean.times" ;
		mean_time:dpl_py_type = "python_datetime" ;
	double time_offset(time) ;
		time_offset:long_name = "Time offset from time_coverage_start" ;
		time_offset:description = "same times as \"First time in record\" " ;
		time_offset:units = "seconds since 2006-10-23 18:19:59 UTC" ;
		time_offset:dpl_py_binding = "dne" ;
	short start_time(time, time_vector) ;
		start_time:long_name = "First Time in record" ;
		start_time:description = "time of first laser shot in averaging interval" ;
		start_time:dpl_py_binding = "dne" ;
	float range_resolution ;
		range_resolution:long_name = "Range resolution" ;
		range_resolution:description = "vertical distance between data points after averaging" ;
		range_resolution:units = "meters" ;
		range_resolution:dpl_py_binding = "dne" ;
	float time_average ;
		time_average:long_name = "Time Averaging Width" ;
		time_average:description = "Time between data points after averaging" ;
		time_average:units = "seconds" ;
		time_average:dpl_py_binding = "dne" ;
	float range(range) ;
		range:standard_name = "projection_range_coodinate" ;
		range:long_name = "range_to_measurement_volume" ;
		range:units = "meters" ;
		range:spacing_is_constant = "yes" ;
		range:meters_to_center_of_first_gate = 0.0 ; // FIXME in netcdf generation
		range:axis = "radial_range_coodinate" ;
		range:dpl_py_binding = "rs_mean.msl_altitudes" ;
	double latitude(time) ;
                latitude:standard_name = "latitude" ;
                latitude:units = "degrees_north" ;
		latitude:dpl_py_binding = "rs_mean.latitude" ;
        double longitude(time) ;
                longitude:standard_name = "longitude" ;
                longitude:units = "degrees_east" ;
		longitude:dpl_py_binding = "rs_mean.longitude" ;
        double altitude(time) ;
                altitude:standard_name = "altitude" ;
                altitude:units = "meters" ;
                altitude:positive = "up" ;
		altitude:dpl_py_binding = "rs_mean.GPS_MSL_Alt" ;
        double telescope_roll_angle_offset(time) ;
                telescope_roll_angle_offset:long_name = "Telescope Mounting Roll Angle Offset" ;
                telescope_roll_angle_offset:description = "Telescope Mount Roll Angle Relative to aircraft up measured clockwise" ;
                telescope_roll_angle_offset:units = "degrees" ;
                		telescope_roll_angle_offset:range = -180.0, 360.0 ;
				telescope_roll_angle_offset:dpl_py_binding = "rs_mean.telescope_roll_angle_offset" ;

        double roll(time) ;
                roll:standard_name = "roll" ;
                roll:units = "degrees" ;
                roll:positive = "left side up looking forward" ;
		roll:dpl_py_binding = "rs_mean.roll_angle" ;

        double pitch(time) ;
                pitch:standard_name = "pitch" ;
                pitch:units = "degrees" ;
                pitch:positive = "up at front" ;
		pitch:dpl_py_binding = "rs_mean.pitch_angle" ;

        double heading(time) ;
                heading:standard_name = "heading" ;
                heading:units = "degrees_true" ;
		heading:dpl_py_binding = "rs_mean.heading" ;
        double drift(time) ;
                drift:standard_name = "drift" ;
                drift:units = "degrees" ;
		drift:dpl_py_binding = "rs_mean.drift" ;
		
	float aeri_btemp_wavenumber(aeri_btemp_wavenumber) ;
		aeri_btemp_wavenumber:long_name = "Wave number" ;
		aeri_btemp_wavenumber:units = "cm^-1" ;
		aeri_btemp_wavenumber:missing_value = 9.96920996838687e+36 ;
		aeri_btemp_wavenumber:dpl_py_binding = "dne" ;
	float aeri_btemp(time, aeri_btemp_wavenumber) ;
		aeri_btemp:long_name = "AERI Brightness Temperature" ;
		aeri_btemp:units = "degK" ;
		aeri_btemp:missing_value = 9.96920996838687e+36 ;
		aeri_btemp:dpl_py_binding = "dne" ;
	float mwr_watervapor(time) ;
		mwr_watervapor:long_name = "MWR Water vapor along LOS path" ;
		mwr_watervapor:units = "cm" ;
		mwr_watervapor:missing_value = 9.96920996838687e+36 ;
		mwr_watervapor:dpl_py_binding = "dne" ;
	float mwr_liquidwater(time) ;
		mwr_liquidwater:long_name = "MWR Liquid water along LOS path" ;
		mwr_liquidwater:units = "g/m^2" ;
		mwr_liquidwater:missing_value = 9.96920996838687e+36 ;
		mwr_liquidwater:dpl_py_binding = "dne" ;
	float aeri_mean_rad_wavenumber_ch1(aeri_mean_rad_wavenumber_ch1) ;
		aeri_mean_rad_wavenumber_ch1:long_name = "Wave number" ;
		aeri_mean_rad_wavenumber_ch1:units = "cm^-1" ;
		aeri_mean_rad_wavenumber_ch1:missing_value = 9.96920996838687e+36 ;
		aeri_mean_rad_wavenumber_ch1:dpl_py_binding = "dne" ;
	float aeri1_mean_rad(time, aeri_mean_rad_wavenumber_ch1) ;
		aeri1_mean_rad:long_name = "Downwelling radiance interpolated to standard wavenumber scale Channel 1" ;
		aeri1_mean_rad:units = "mw/(m2 sr cm-1)" ;
		aeri1_mean_rad:missing_value = 9.96920996838687e+36 ;
		aeri1_mean_rad:dpl_py_binding = "dne" ;
	int aeri_qc(time) ;
		aeri_qc:long_name = "Aeri Quality" ;
		aeri_qc:bit_0 = "channel 1" ;
		aeri_qc:bit_1 = "channel 2" ;
		aeri_qc:missing_value = -1 ;
		aeri_qc:dpl_py_binding = "dne" ;
	float aeri_mean_rad_wavenumber_ch2(aeri_mean_rad_wavenumber_ch2) ;
		aeri_mean_rad_wavenumber_ch2:long_name = "Wave number" ;
		aeri_mean_rad_wavenumber_ch2:units = "cm^-1" ;
		aeri_mean_rad_wavenumber_ch2:missing_value = 9.96920996838687e+36 ;
		aeri_mean_rad_wavenumber_ch2:dpl_py_binding = "dne" ;
	float aeri2_mean_rad(time, aeri_mean_rad_wavenumber_ch2) ;
		aeri2_mean_rad:long_name = "Downwelling radiance interpolated to standard wavenumber scale Channel 2" ;
		aeri2_mean_rad:units = "mw/(m2 sr cm-1)" ;
		aeri2_mean_rad:missing_value = 9.96920996838687e+36 ;
		aeri2_mean_rad:dpl_py_binding = "dne" ;
	float aeri1_pca_mean_rad(time, aeri_mean_rad_wavenumber_ch1) ;
		aeri1_pca_mean_rad:long_name = "PCA Filtered Downwelling radiance interpolated to standard wavenumber scale Channel 1" ;
		aeri1_pca_mean_rad:units = "mw/(m2 sr cm-1)" ;
		aeri1_pca_mean_rad:missing_value = 9.96920996838687e+36 ;
		aeri1_pca_mean_rad:dpl_py_binding = "dne" ;
	float aeri2_pca_mean_rad(time, aeri_mean_rad_wavenumber_ch2) ;
		aeri2_pca_mean_rad:long_name = "PCA Filtered Downwelling radiance interpolated to standard wavenumber scale Channel 2" ;
		aeri2_pca_mean_rad:units = "mw/(m2 sr cm-1)" ;
		aeri2_pca_mean_rad:missing_value = 9.96920996838687e+36 ;
		aeri2_pca_mean_rad:dpl_py_binding = "dne" ;
	float beta_m(calibration, range) ;
		beta_m:long_name = "Raob molecular scattering cross section per unit volume" ;
		beta_m:units = "1/meter" ;
		beta_m:plot_scale = "logarithmic" ;
		beta_m:dpl_py_binding = "rs_Cxx.beta_r" ;
	float transmitted_energy(time) ;
		transmitted_energy:long_name = "Transmitted Energy" ;
		transmitted_energy:units = "Joules" ;
		transmitted_energy:missing_value = 9.96920996838687e+36 ;
		transmitted_energy:dpl_py_binding = "rs_mean.transmitted_energy" ;
	float piezovoltage(time) ;
		piezovoltage:long_name = "piezovoltage" ;
		piezovoltage:units = "Volts" ;
		piezovoltage:missing_value = 9.96920996838687e+36 ;
		piezovoltage:dpl_py_binding = "dne" ;
	int num_seeded_shots(time) ;
		num_seeded_shots:long_name = "Number of Seeded Shots" ;
		num_seeded_shots:missing_value = -1 ;
		num_seeded_shots:dpl_py_binding = "rs_mean.seeded_shots" ;
	int num_shots(time) ;
		num_shots:long_name = "Number of Shots" ;
		num_shots:missing_value = -1 ;
		num_shots:dpl_py_binding = "rs_mean.shot_count" ;
	float seed_quality(time) ;
		seed_quality:long_name = "Laser Seeding Quality" ;
		seed_quality:description = "The ratio of seeded shots to total shots. Only seeded shot data is stored and processed.  A low seed ratio can result in low noise resistance." ;
		seed_quality:missing_value = 9.96920996838687e+36 ;
		seed_quality:range = 0., 1. ;
		seed_quality:dpl_py_binding = "dne" ;
	float frequency_quality(time) ;
		frequency_quality:long_name = "Laser Frequency Quality" ;
		frequency_quality:description = "An ratio average of how good the frequency lock is per raw interval. A low value can result in poor separation of molecular and aerosol counts." ;
		frequency_quality:missing_value = 9.96920996838687e+36 ;
		frequency_quality:range = 0., 1. ;
		frequency_quality:dpl_py_binding = "dne" ;
	float lock_quality(time) ;
		lock_quality:long_name = "Laser Lock Quality" ;
		lock_quality:description = "A ratio of likely locked intervals (frequency_quality>=.5) to seeded intervals.  A low value can result in poor separation of molecular and aerosol counts." ;
		lock_quality:missing_value = 9.96920996838687e+36 ;
		lock_quality:range = 0., 1. ;
		lock_quality:dpl_py_binding = "dne" ;
	float mol_cal_pulse(time) ;
		mol_cal_pulse:long_name = "Molecular calibration pulse" ;
		mol_cal_pulse:description = "Sum of photon counts in the molecular channel due to light scattered with the telescope." ;
		mol_cal_pulse:units = "counts" ;
		mol_cal_pulse:missing_value = 9.96920996838687e+36 ;
		mol_cal_pulse:dpl_py_binding = "rs_mean.molecular_cal_pulse" ;
	float c_pol_dark_count(time) ;
		c_pol_dark_count:long_name = "Cross Polarization Dark Count FIXME dark counts need alt" ;
		c_pol_dark_count:description = "total counts per averaging interval(eg. one range, one time)" ;
		c_pol_dark_count:units = "counts" ;
		c_pol_dark_count:missing_value = 9.96920996838687e+36 ;
		c_pol_dark_count:dpl_py_binding = "rs_mean.c_pol_dark_counts" ;
	float mol_dark_count(time) ;
		mol_dark_count:long_name = "Molecular Dark Count" ;
		mol_dark_count:description = "total counts per averaging interval(eg. one range, one time)" ;
		mol_dark_count:units = "counts" ;
		mol_dark_count:missing_value = 9.96920996838687e+36 ;
		mol_dark_count:dpl_py_binding = "rs_mean.mol_dark_counts" ;
	float combined_dark_count_lo(time) ;
		combined_dark_count_lo:long_name = "Low Gain Combined Dark Count" ;
		combined_dark_count_lo:description = "total counts per averaging interval(eg. one range, one time)" ;
		combined_dark_count_lo:units = "counts" ;
		combined_dark_count_lo:missing_value = 9.96920996838687e+36 ;
		combined_dark_count_lo:dpl_py_binding = "rs_mean.c_lo_dark_counts" ;
	float combined_dark_count_hi(time) ;
		combined_dark_count_hi:long_name = "High Gain Combined Dark Count" ;
		combined_dark_count_hi:description = "total counts per averaging interval(eg. one range, one time)" ;
		combined_dark_count_hi:units = "counts" ;
		combined_dark_count_hi:missing_value = 9.96920996838687e+36 ;
		combined_dark_count_hi:dpl_py_binding = "rs_mean.c_hi_dark_counts" ;
	float combined_gain(calibration) ;
		combined_gain:long_name = "Combined Gain Factor" ;
		combined_gain:description = "Low Gain level * Factor ~ High Gain level" ;
		combined_gain:dpl_py_binding = "rs_constants.hi_to_low_combined_channel_gain_ratio" ;
	float combined_merge_threshhold(calibration) ;
		combined_merge_threshhold:long_name = "Combined Merge Threshhold" ;
		combined_merge_threshhold:dpl_py_binding = "rs_constants.combined_channel_merge_threshhold" ;
	float polarization_cross_talk(calibration) ;
		polarization_cross_talk:long_name = "Polarization Cross Talk" ;
		polarization_cross_talk:dpl_py_binding = "rs_constants.polarization_cross_talk" ;
	float wfov_to_combined_gain_ratio(calibration) ;
		wfov_to_combined_gain_ratio:long_name = "WFOV to Combined Gain" ;
		wfov_to_combined_gain_ratio:dpl_py_binding = "rs_constants.wfov_to_combined_gain_ratio" ;
	float combined_to_cross_pol_gain_ratio(calibration) ;
		combined_to_cross_pol_gain_ratio:long_name = "Combined to Cross Pol Gain" ;
		combined_to_cross_pol_gain_ratio:dpl_py_binding = "rs_constants.combined_to_cross_pol_gain_ratio" ;
	float molecular_to_wfov_gain_ratio(calibration) ;
		molecular_to_wfov_gain_ratio:long_name = "Molecular to WFOV Gain" ;
		molecular_to_wfov_gain_ratio:dpl_py_binding = "rs_constants.molecular_to_wfov_gain_ratio" ;
	float geo_cor(calibration, bin_range) ;
		geo_cor:long_name = "Overlap correction" ;
		geo_cor:description = "Geometric overlap correction in raw range bins" ;
		geo_cor:units = " " ;
		geo_cor:missing_value = 9.96920996838687e+36 ;
		geo_cor:plot_scale = "logarithmic" ;
		geo_cor:dpl_py_binding = "geo_corr" ;
	int od_norm_index ;
		od_norm_index:long_name = "Optical depth normalization index FIXME shouldn't be needed" ;
		od_norm_index:dpl_py_binding = "rs_inv.od_norm_index" ;
	float od(time, range) ;
		od:long_name = "Aerosol + Molecular Optical Depth" ;
		od:units = " " ;
		od:missing_value = 9.96920996838687e+36 ;
		od:insufficient_data = 9.96920996838687e+36 ;
		od:plot_scale = "logarithmic" ;
		od:dpl_py_binding = "rs_inv.optical_depth" ;
	float profile_od(profile_time,range) ;
		profile_od:long_name = "Aerosol + Molecular Optical Depth Profile" ;
		profile_od:units = " " ;
		profile_od:missing_value = 9.96920996838687e+36 ;
		profile_od:insufficient_data = 9.96920996838687e+36 ;
		profile_od:plot_scale = "logarithmic" ;
		profile_od:dpl_py_binding = "profiles.inv.optical_depth" ;
	float profile_extinction(profile_time,range) ;
		profile_extinction:long_name = "Aerosol + Molecular Extinction Profile" ;
		profile_extinction:units = " " ;
		profile_extinction:missing_value = 9.96920996838687e+36 ;
		profile_extinction:insufficient_data = 9.96920996838687e+36 ;
		profile_extinction:plot_scale = "logarithmic" ;
		profile_extinction:dpl_py_binding = "profiles.inv.extinction" ;
	float extinction(time,range) ;
		extinction:long_name = "Aerosol + Molecular Extinction Profile" ;
		extinction:units = " " ;
		extinction:missing_value = 9.96920996838687e+36 ;
		extinction:insufficient_data = 9.96920996838687e+36 ;
		extinction:plot_scale = "logarithmic" ;
		extinction:dpl_py_binding = "rs_inv.extinction" ;
	float od_aerosol(time, range) ;
		od_aerosol:long_name = "Aerosol Optical Depth" ;
		od_aerosol:units = " " ;
		od_aerosol:missing_value = 9.96920996838687e+36 ;
		od_aerosol:insufficient_data = 9.96920996838687e+36 ;
		od_aerosol:plot_scale = "logarithmic" ;
		od_aerosol:dpl_py_binding = "rs_inv.optical_depth_aerosol" ;
	float profile_od_aerosol(profile_time,range) ;
		profile_od_aerosol:long_name = "Aerosol Optical Depth Profile" ;
		profile_od_aerosol:units = " " ;
		profile_od_aerosol:missing_value = 9.96920996838687e+36 ;
		profile_od_aerosol:insufficient_data = 9.96920996838687e+36 ;
		profile_od_aerosol:plot_scale = "logarithmic" ;
		profile_od_aerosol:dpl_py_binding = "profiles.inv.optical_depth_aerosol" ;
	float profile_extinction_aerosol(profile_time,range) ;
		profile_extinction_aerosol:long_name = "Aerosol Extinction Profile" ;
		profile_extinction_aerosol:units = " " ;
		profile_extinction_aerosol:missing_value = 9.96920996838687e+36 ;
		profile_extinction_aerosol:insufficient_data = 9.96920996838687e+36 ;
		profile_extinction_aerosol:plot_scale = "logarithmic" ;
		profile_extinction_aerosol:dpl_py_binding = "profiles.inv.extinction_aerosol" ;
	float extinction_aerosol(time,range) ;
		extinction_aerosol:long_name = "Aerosol Extinction" ;
		extinction_aerosol:units = " " ;
		extinction_aerosol:missing_value = 9.96920996838687e+36 ;
		extinction_aerosol:insufficient_data = 9.96920996838687e+36 ;
		extinction_aerosol:plot_scale = "logarithmic" ;
		extinction_aerosol:dpl_py_binding = "rs_inv.extinction_aerosol" ;
	float radar_backscattercrosssection(time, range) ;
		radar_backscattercrosssection:long_name = "MMCR Backscatter Cross Section" ;
		radar_backscattercrosssection:units = "1/(m sr)" ;
		radar_backscattercrosssection:missing_value = 9.96920996838687e+36 ;
		radar_backscattercrosssection:dpl_py_binding = "dne" ;
	float radar_reflectivity(time, range) ;
		radar_reflectivity:long_name = "MMCR Reflectivity" ;
		radar_reflectivity:units = "dBz" ;
		radar_reflectivity:missing_value = 9.96920996838687e+36 ;
		radar_reflectivity:dpl_py_binding = "dne" ;
	float radar_spectralwidth(time, range) ;
		radar_spectralwidth:long_name = "MMCR Spectral Width" ;
		radar_spectralwidth:units = "m/s" ;
		radar_spectralwidth:missing_value = 9.96920996838687e+36 ;
		radar_spectralwidth:dpl_py_binding = "dne" ;
	float radar_dopplervelocity(time, range) ;
		radar_dopplervelocity:long_name = "MMCR doppler Velocity" ;
		radar_dopplervelocity:units = "m/s" ;
		radar_dopplervelocity:missing_value = 9.96920996838687e+36 ;
		radar_dopplervelocity:dpl_py_binding = "dne" ;
	float effective_diameter_prime(time, range) ;
		effective_diameter_prime:long_name = "lidar/radar effective particle diameter" ;
		effective_diameter_prime:units = "microns" ;
		effective_diameter_prime:description = "Effective diameter directly from the ratio of Lidar Backscatter and Radar Reflectivity; (<volume^2>/<area>)^.25, see Donovan JGR Nov 2001" ;
		effective_diameter_prime:missing_value = 9.96920996838687e+36 ;
		effective_diameter_prime:dpl_py_binding = "dne" ;
	float effective_diameter(time, range) ;
		effective_diameter:long_name = "Effective particle diameter" ;
		effective_diameter:units = "microns" ;
		effective_diameter:description = "Effective particle diameter derived from ratio of Lidar Backscatter and Radar Reflectivity; assuming a gamma size distribution" ;
		effective_diameter:missing_value = 9.96920996838687e+36 ;
		effective_diameter:dpl_py_binding = "dne" ;
	float num_particles(time, range) ;
		num_particles:long_name = "Number density of particles" ;
		num_particles:units = "1/liter" ;
		num_particles:description = "Number of particles per liter derived from ratio of lidar backscatter and radar reflectivity; assuming a gamma size distribution" ;
		num_particles:missing_value = 9.96920996838687e+36 ;
		num_particles:dpl_py_binding = "dne" ;
	float mean_diameter(time, range) ;
		mean_diameter:long_name = "Mean diameter of particles" ;
		mean_diameter:units = "microns" ;
		mean_diameter:description = "Mean diameter of particles derived from the effective diameter and the gamma size distribution" ;
		mean_diameter:missing_value = 9.96920996838687e+36 ;
		mean_diameter:dpl_py_binding = "dne" ;
	float LWC(time, range) ;
		LWC:long_name = "Liquid water content" ;
		LWC:units = "gr/m^3" ;
		LWC:description = "Liquid water content derived from ratio of lidar backscatter and radar reflectivity; assuming a gamma size distribution" ;
		LWC:missing_value = 9.96920996838687e+36 ;
		LWC:dpl_py_binding = "dne" ;
	float beta_a(time, range) ;
		beta_a:long_name = "Particulate extinction cross section per unit volume" ;
		beta_a:units = "1/m" ;
		beta_a:missing_value = 9.96920996838687e+36 ;
		beta_a:plot_scale = "logarithmic" ;
		beta_a:dpl_py_binding = "dne" ;
	float atten_beta_r_backscat(time, range) ;
		atten_beta_r_backscat:long_name = "Attenuated Molecular return" ;
		atten_beta_r_backscat:units = "1/(m sr)" ;
		atten_beta_r_backscat:missing_value = 9.96920996838687e+36 ;
		atten_beta_r_backscat:plot_scale = "logarithmic" ;
		atten_beta_r_backscat:dpl_py_binding = "rs_inv.atten_beta_a_backscat" ;
	float profile_atten_beta_r_backscat(range) ;
		profile_atten_beta_r_backscat:long_name = "Attenuated Molecular Profile" ;
		profile_atten_beta_r_backscat:units = "1/(m sr)" ;
		profile_atten_beta_r_backscat:missing_value = 9.96920996838687e+36 ;
		profile_atten_beta_r_backscat:plot_scale = "logarithmic" ;
		profile_atten_beta_r_backscat:dpl_py_binding = "profiles.inv.atten_beta_a_backscat" ;
	float circular_depol(time, range) ;
		circular_depol:long_name = "Circular depolarization ratio for particulate" ;
		circular_depol:description = "left circular return divided by right circular return" ;
		circular_depol:units = " " ;
		circular_depol:missing_value = 9.96920996838687e+36 ;
		circular_depol:plot_scale = "logarithmic" ;
		circular_depol:dpl_py_binding = "rs_inv.circular_depol" ;
	float linear_depol(time, range) ;
		linear_depol:long_name = "Linear depolarization ratio for particulate" ;
		linear_depol:description = "Linear depolarization return" ;
		linear_depol:units = " " ;
		linear_depol:missing_value = 9.96920996838687e+36 ;
		linear_depol:plot_scale = "logarithmic" ;
		linear_depol:dpl_py_binding = "rs_inv.linear_depol" ;
	float profile_circular_depol(profile_time,range) ;
		profile_circular_depol:long_name = "Circular depolarization ratio profile for particulate" ;
		profile_circular_depol:description = "left circular return divided by right circular return" ;
		profile_circular_depol:units = " " ;
		profile_circular_depol:missing_value = 9.96920996838687e+36 ;
		profile_circular_depol:plot_scale = "logarithmic" ;
		profile_circular_depol:dpl_py_binding = "profiles.inv.circular_depol" ;
	float profile_linear_depol(profile_time,range) ;
		profile_linear_depol:long_name = "Linear depolarization ratio profile for particulate" ;
		profile_linear_depol:description = "??? return" ;
		profile_linear_depol:units = " " ;
		profile_linear_depol:missing_value = 9.96920996838687e+36 ;
		profile_linear_depol:plot_scale = "logarithmic" ;
		profile_linear_depol:dpl_py_binding = "profiles.inv.linear_depol" ;
	float beta_a_backscat_parallel(time, range) ;
		beta_a_backscat_parallel:long_name = "Particulate nondepolarized backscatter cross section per unit volume" ;
		beta_a_backscat_parallel:units = "1/(m sr)" ;
		beta_a_backscat_parallel:missing_value = 9.96920996838687e+36 ;
		beta_a_backscat_parallel:plot_scale = "logarithmic" ;
		beta_a_backscat_parallel:dpl_py_binding = "rs_inv.beta_a_backscat_par" ;
	float profile_beta_a_backscat_parallel(profile_time,range) ;
		profile_beta_a_backscat_parallel:long_name = "Particulate nondepolarized backscatter cross section profile" ;
		profile_beta_a_backscat_parallel:units = "1/(m sr)" ;
		profile_beta_a_backscat_parallel:missing_value = 9.96920996838687e+36 ;
		profile_beta_a_backscat_parallel:plot_scale = "logarithmic" ;
		profile_beta_a_backscat_parallel:dpl_py_binding = "profiles.inv.beta_a_backscat_par" ;
	float beta_a_backscat_perpendicular(time, range) ;
		beta_a_backscat_perpendicular:long_name = "Particulate depolarized backscatter cross section per unit volume" ;
		beta_a_backscat_perpendicular:units = "1/(m sr)" ;
		beta_a_backscat_perpendicular:missing_value = 9.96920996838687e+36 ;
		beta_a_backscat_perpendicular:plot_scale = "logarithmic" ;
		beta_a_backscat_perpendicular:dpl_py_binding = "rs_inv.beta_a_backscat_perp" ;
	float profile_beta_a_backscat_perpendicular(profile_time,range) ;
		profile_beta_a_backscat_perpendicular:long_name = "Particulate depolarized backscatter cross section profile" ;
		profile_beta_a_backscat_perpendicular:units = "1/(m sr)" ;
		profile_beta_a_backscat_perpendicular:missing_value = 9.96920996838687e+36 ;
		profile_beta_a_backscat_perpendicular:plot_scale = "logarithmic" ;
		profile_beta_a_backscat_perpendicular:dpl_py_binding = "profiles.inv.beta_a_backscat_perp" ;
	float beta_a_backscat(time, range) ;
		beta_a_backscat:long_name = "Particulate backscatter cross section per unit volume" ;
		beta_a_backscat:units = "1/(m sr)" ;
		beta_a_backscat:missing_value = 9.96920996838687e+36 ;
		beta_a_backscat:plot_scale = "logarithmic" ;
		beta_a_backscat:dpl_py_binding = "rs_inv.beta_a_backscat" ;
	float profile_beta_a_backscat(profile_time,range) ;
		profile_beta_a_backscat:long_name = "Particulate backscatter cross section profile" ;
		profile_beta_a_backscat:units = "1/(m sr)" ;
		profile_beta_a_backscat:missing_value = 9.96920996838687e+36 ;
		profile_beta_a_backscat:plot_scale = "logarithmic" ;
		profile_beta_a_backscat:dpl_py_binding = "profiles.inv.beta_a_backscat" ;
	float Na(time, range) ;
		Na:long_name = "Inverted Aerosol" ;
		Na:units = " " ;
		Na:dpl_py_binding = "rs_inv.Na" ;
	float Nm(time, range) ;
		Nm:long_name = "Inverted Molecular" ;
		Nm:units = " " ;
		Nm:dpl_py_binding = "rs_inv.Nm" ;
	float Ncp(time, range) ;
		Ncp:long_name = "Inverted Cross Polarization" ;
		Ncp:units = " " ;
		Ncp:dpl_py_binding = "rs_inv.Ncp" ;
	float profile_Na(profile_time,range) ;
		profile_Na:long_name = "Inverted Aerosol Profile" ;
		profile_Na:units = " " ;
		profile_Na:dpl_py_binding = "profiles.inv.Na" ;
	float profile_Nm(profile_time,range) ;
		profile_Nm:long_name = "Inverted Molecular Profile" ;
		profile_Nm:units = " " ;
		profile_Nm:dpl_py_binding = "profiles.inv.Nm" ;
	float profile_Ncp(profile_time,range) ;
		profile_Ncp:long_name = "Inverted Cross Polarization Profile" ;
		profile_Ncp:units = " " ;
		profile_Ncp:dpl_py_binding = "profiles.inv.Ncp" ;

	int qc_mask(time, range) ;
		qc_mask:long_name = "Quality Mask" ;
		qc_mask:description = "Quality mask bitfield.  Unused bits are always high" ;
		qc_mask:missing_value = 0 ;
		qc_mask:_Unsigned = "true" ;
		qc_mask:bit_0 = "complete_mask" ;
		qc_mask:bit_0_description = "data is good.  and of bits 1-9" ;
		qc_mask:bit_1 = "lidar_ok_mask" ;
		qc_mask:bit_1_description = "lidar data is present" ;
		qc_mask:bit_2 = "lock_quality_mask" ;
		qc_mask:bit_2_description = "laser is locked to iodine filter wavelength" ;
		qc_mask:bit_3 = "seed_quality_mask" ;
		qc_mask:bit_3_description = "laser wavelength is locked to seed laser" ;
		qc_mask:bit_4 = "mol_count_snr_mask" ;
		qc_mask:bit_4_description = "molecular signal/photon counting error in molecular signal is above specified threshhold" ;
		qc_mask:bit_5 = "backscat_snr_mask" ;
		qc_mask:bit_5_description = "backscatter cross-section/photon counting error in backscatter cross-section is above specified threshhold" ;
		qc_mask:bit_6 = "mol_lost_mask" ;
		qc_mask:bit_6_description = "number of molecular photon counts is above specified threshhold" ;
		qc_mask:bit_7 = "min_backscat_mask" ;
		qc_mask:bit_7_description = "lidar backscatter cross-section is above specified threshhold" ;
		qc_mask:bit_8 = "radar_backscat_mask" ;
		qc_mask:bit_8_description = "radar backscatter cross-section is above specified threshhold" ;
		qc_mask:bit_9 = "radar_ok_mask" ;
		qc_mask:bit_9_description = "radar data is present" ;
		qc_mask:bit_10 = "aeri_ok_mask" ;
		qc_mask:bit_10_description = "aeri data is present" ;
		qc_mask:bit_11 = "aeri_qc_mask" ;
		qc_mask:bit_11_description = "aeri data has passed a quality check" ;
		qc_mask:dpl_py_binding = "rs_inv.qc_mask" ;
	float std_beta_a_backscat(time, range) ;
		std_beta_a_backscat:long_name = "Std dev of backscat cross section (photon counting)" ;
		std_beta_a_backscat:units = "1/(m sr)" ;
		std_beta_a_backscat:missing_value = 9.96920996838687e+36 ;
		std_beta_a_backscat:plot_scale = "logarithmic" ;
		std_beta_a_backscat:dpl_py_binding = "rs_inv.std_beta_a_backscat" ;
	float mwr_frequency(mwr_frequency) ;
		mwr_frequency:long_name = "Frequency" ;
		mwr_frequency:units = "GHz" ;
		mwr_frequency:missing_value = 9.96920996838687e+36 ;
		mwr_frequency:dpl_py_binding = "dne" ;
	float mwr_btemp(time, mwr_frequency) ;
		mwr_btemp:long_name = "MWR Brightness Temperature" ;
		mwr_btemp:units = "degK" ;
		mwr_btemp:missing_value = 9.96920996838687e+36 ;
		mwr_btemp:dpl_py_binding = "dne" ;

	int sweep_number(sweep) ;
                sweep_number:standard_name = "sweep_index_number_0_based" ;
                sweep_number:_FillValue = -9999 ;

        char sweep_mode(sweep, string_length_short) ;
                sweep_mode:standard_name = "scan_mode_for_sweep" ;
                sweep_mode:options = "sector, coplane, rhi, vertical_pointing, idle, azimuth_surveillance, elevation_surveillance, sunscan, pointing, calibration, manual_ppi, manual_rhi" ;

        float fixed_angle(sweep) ;
                fixed_angle:standard_name = "beam_target_fixed_angle" ;
                fixed_angle:units = "degrees" ;
                fixed_angle:_FillValue = -9999.f ;

        int sweep_start_ray_index(sweep) ;
                sweep_start_ray_index:standard_name = "index_of_first_ray_in_sweep" ;
                sweep_start_ray_index:_FillValue = -9999 ;
        int sweep_end_ray_index(sweep) ;
                sweep_end_ray_index:standard_name = "index_of_last_ray_in_sweep" ;
                sweep_end_ray_index:_FillValue = -9999 ;

// global attributes:
                :dpl_py_template = "hsrl_cfradial.cdl" ;
                :dpl_py_template_version = 20120526 ;
		:time_zone = "UTC" ;
	        :Conventions = "CF/Radial instrument_parameters" ;
                :version = "1.2" ;
		:title = "GV HSRL lidar data";
		:institution = "EOL/NCAR" ;
		:references = "eol_hsrl_python" ;
		:source = "GV HSRL" ;
		:instrument_name = "GV HSRL" ;
		:comment = "" ;
		:history = "" ;
		:platform_is_mobile = "true" ;
}
