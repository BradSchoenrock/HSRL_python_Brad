netcdf out {
dimensions:
	raw_time = UNLIMITED ;
	bin_range = 0 ;
	profile_time = 1;
	time_vector = 8 ;
variables:
	int base_time ;
		base_time:string = "2006-10-23 18:19:59 UTC" ;
		base_time:long_name = "Base seconds since Unix Epoch" ;
		base_time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		base_time:dpl_py_binding = "dne" ;
	double raw_time(raw_time) ;
		raw_time:long_name = "Raw Time" ;
		raw_time:units = "seconds since 2006-10-23 18:19:59 UTC" ;
		raw_time:dpl_py_binding = "rs_raw.times" ;
		raw_time:dpl_py_type = "python_datetime" ;
	float altitude(bin_range) ;
		altitude:long_name = "Height above lidar" ;
		altitude:units = "meters" ;
		altitude:dpl_py_binding = "rs_raw.msl_altitudes" ;
	float transmitted_energy(raw_time) ;
		transmitted_energy:long_name = "Transmitted Energy" ;
		transmitted_energy:units = "Joules" ;
		transmitted_energy:dpl_py_binding = "rs_raw.transmitted_energy" ;
	float transmitted_1064_energy(raw_time) ;
		transmitted_1064_energy:long_name = "Transmitted 1064 IR Energy" ;
		transmitted_1064_energy:units = "Joules" ;
		transmitted_1064_energy:dpl_py_binding = "rs_raw.transmitted_1064_energy" ;
	int num_seeded_shots(raw_time) ;
		num_seeded_shots:long_name = "Number of Seeded Shots" ;
		num_seeded_shots:missing_value = -1 ;
		num_seeded_shots:dpl_py_binding = "rs_raw.seeded_shots" ;
	int num_shots(raw_time) ;
		num_shots:long_name = "Number of Shots" ;
		num_shots:missing_value = -1 ;
		num_shots:dpl_py_binding = "rs_raw.shot_count" ;
	float mol_cal_pulse(raw_time) ;
		mol_cal_pulse:long_name = "Molecular calibration pulse" ;
		mol_cal_pulse:description = "Sum of photon counts in the molecular channel due to light scattered with the telescope." ;
		mol_cal_pulse:units = "counts" ;
		mol_cal_pulse:dpl_py_binding = "rs_raw.molecular_cal_pulse" ;
	int molecular_counts(raw_time, bin_range) ;
		molecular_counts:long_name = "Molecular Photon Counts" ;
		molecular_counts:description = "Raw counts, per averaging interval with pileup applied" ;
		molecular_counts:units = "counts" ;
		molecular_counts:missing_value = -1 ;
		molecular_counts:plot_scale = "logarithmic" ;
		molecular_counts:dpl_py_binding = "rs_raw.molecular_counts" ;
	int molecular_i2a_counts(raw_time, bin_range) ;
		molecular_i2a_counts:long_name = "Molecular I2A Photon Counts" ;
		molecular_i2a_counts:description = "Raw counts, per averaging interval with pileup applied" ;
		molecular_i2a_counts:units = "counts" ;
		molecular_i2a_counts:missing_value = -1 ;
		molecular_i2a_counts:plot_scale = "logarithmic" ;
		molecular_i2a_counts:dpl_py_binding = "rs_raw.molecular_i2a_counts" ;
	int molecular_wfov_counts(raw_time, bin_range) ;
		molecular_wfov_counts:long_name = "Molecular WFOV Photon Counts" ;
		molecular_wfov_counts:description = "Raw counts, per averaging interval with pileup applied" ;
		molecular_wfov_counts:units = "counts" ;
		molecular_wfov_counts:missing_value = -1 ;
		molecular_wfov_counts:plot_scale = "logarithmic" ;
		molecular_wfov_counts:dpl_py_binding = "rs_raw.molecular_wfov_counts" ;
	int combined_counts_lo(raw_time, bin_range) ;
		combined_counts_lo:long_name = "Low Gain Combined Photon Counts" ;
		combined_counts_lo:description = "Raw counts, per averaging interval with pileup applied" ;
		combined_counts_lo:units = "counts" ;
		combined_counts_lo:missing_value = -1 ;
		combined_counts_lo:plot_scale = "logarithmic" ;
		combined_counts_lo:dpl_py_binding = "rs_raw.combined_lo_counts" ;
	int combined_counts_hi(raw_time, bin_range) ;
		combined_counts_hi:long_name = "High Gain Combined Photon Counts" ;
		combined_counts_hi:description = "Raw counts, per averaging interval with pileup applied" ;
		combined_counts_hi:units = "counts" ;
		combined_counts_hi:missing_value = -1 ;
		combined_counts_hi:plot_scale = "logarithmic" ;
		combined_counts_hi:dpl_py_binding = "rs_raw.combined_hi_counts" ;
	int combined_counts(raw_time, bin_range) ;
		combined_counts:long_name = "Combined Photon Counts" ;
		combined_counts:description = "Raw counts, per averaging interval with pileup applied" ;
		combined_counts:units = "counts" ;
		combined_counts:missing_value = -1 ;
		combined_counts:plot_scale = "logarithmic" ;
		combined_counts:dpl_py_binding = "rs_raw.combined_counts" ;
	int combined_1064_counts(raw_time, bin_range) ;
		combined_1064_counts:long_name = "1064 IR Combined Photon Counts" ;
		combined_1064_counts:description = "Raw counts, per averaging interval with pileup applied" ;
		combined_1064_counts:units = "counts" ;
		combined_1064_counts:missing_value = -1 ;
		combined_1064_counts:plot_scale = "logarithmic" ;
		combined_1064_counts:dpl_py_binding = "rs_raw.combined_1064_counts" ;
	int cross_counts(raw_time, bin_range) ;
		cross_counts:long_name = "Cross Polarized Photon Counts" ;
		cross_counts:description = "Raw counts, per averaging interval with pileup applied" ;
		cross_counts:units = "counts" ;
		cross_counts:missing_value = -1 ;
		cross_counts:plot_scale = "logarithmic" ;
		cross_counts:dpl_py_binding = "rs_raw.cross_pol_counts" ;
	float c_pol_dark_count(raw_time) ;
		c_pol_dark_count:long_name = "Cross Polarization Dark Count" ;
		c_pol_dark_count:description = "total counts per averaging interval(eg. one altitude, one time)" ;
		c_pol_dark_count:units = "counts" ;
		c_pol_dark_count:dpl_py_binding = "rs_raw.c_pol_dark_counts" ;
	float mol_i2a_dark_count(raw_time) ;
		mol_i2a_dark_count:long_name = "Molecular I2A Dark Count" ;
		mol_i2a_dark_count:description = "total counts per averaging interval(eg. one altitude, one time)" ;
		mol_i2a_dark_count:units = "counts" ;
		mol_i2a_dark_count:dpl_py_binding = "rs_raw.mol_i2a_dark_counts" ;
	float mol_dark_count(raw_time) ;
		mol_dark_count:long_name = "Molecular Dark Count" ;
		mol_dark_count:description = "total counts per averaging interval(eg. one altitude, one time)" ;
		mol_dark_count:units = "counts" ;
		mol_dark_count:dpl_py_binding = "rs_raw.mol_dark_counts" ;
	float combined_dark_count_lo(raw_time) ;
		combined_dark_count_lo:long_name = "Low Gain Combined Dark Count" ;
		combined_dark_count_lo:description = "total counts per averaging interval(eg. one altitude, one time)" ;
		combined_dark_count_lo:units = "counts" ;
		combined_dark_count_lo:dpl_py_binding = "rs_raw.c_lo_dark_counts" ;
	float combined_dark_count_hi(raw_time) ;
		combined_dark_count_hi:long_name = "High Gain Combined Dark Count" ;
		combined_dark_count_hi:description = "total counts per averaging interval(eg. one altitude, one time)" ;
		combined_dark_count_hi:units = "counts" ;
		combined_dark_count_hi:dpl_py_binding = "rs_raw.c_hi_dark_counts" ;
	float combined_1064_dark_count(raw_time) ;
		combined_1064_dark_count:long_name = "Combined 1064 Dark Count" ;
		combined_1064_dark_count:description = "total counts per averaging interval(eg. one altitude, one time)" ;
		combined_1064_dark_count:units = "counts" ;
		combined_1064_dark_count:dpl_py_binding = "rs_raw.combined_1064_dark_count" ;
	float combined_dark_count(raw_time) ;
		combined_dark_count:long_name = "Combined Dark Count" ;
		combined_dark_count:description = "total counts per averaging interval(eg. one altitude, one time)" ;
		combined_dark_count:units = "counts" ;
		combined_dark_count:dpl_py_binding = "rs_raw.c_dark_counts" ;

// global attributes:
		:dpl_py_template = "hsrl3_raw.cdl" ;
		:dpl_py_template_version = 20150813 ;
		:time_zone = "UTC" ;
}
