netcdf out {
dimensions:
	altitude = 0 ;
    profile_time = 1;
	time_vector = 8 ;
variables:
	int base_time ;
		base_time:string = "2006-10-23 18:19:59 UTC" ;
		base_time:long_name = "Base seconds since Unix Epoch" ;
		base_time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		base_time:dpl_py_binding = "dne" ;
	short first_time(time_vector) ;
		first_time:long_name = "First Time in file" ;
		first_time:dpl_py_binding = "dne" ;
	short last_time(time_vector) ;
		last_time:long_name = "Last Time in file" ;
		last_time:dpl_py_binding = "dne" ;
	float altitude(altitude) ;
		altitude:long_name = "Height above lidar" ;
		altitude:units = "meters" ;
		altitude:dpl_py_binding = "rs_mean.msl_altitudes" ;
	float profile_od(profile_time,altitude) ;
		profile_od:long_name = "Optical depth of particulate Profile" ;
		profile_od:units = " " ;
		profile_od:missing_value = 9.96920996838687e+36 ;
		profile_od:insufficient_data = 9.96920996838687e+36 ;
		profile_od:plot_scale = "logarithmic" ;
		profile_od:dpl_py_binding = "profiles.inv.optical_depth" ;
	float profile_extinction(profile_time,altitude) ;
		profile_extinction:long_name = "Extinction Profile" ;
		profile_extinction:units = " " ;
		profile_extinction:missing_value = 9.96920996838687e+36 ;
		profile_extinction:insufficient_data = 9.96920996838687e+36 ;
		profile_extinction:plot_scale = "logarithmic" ;
		profile_extinction:dpl_py_binding = "profiles.inv.extinction" ;
	float profile_atten_beta_r_backscat(altitude) ;
		profile_atten_beta_r_backscat:long_name = "Attenuated Molecular Profile" ;
		profile_atten_beta_r_backscat:units = "1/(m sr)" ;
		profile_atten_beta_r_backscat:missing_value = 9.96920996838687e+36 ;
		profile_atten_beta_r_backscat:plot_scale = "logarithmic" ;
		profile_atten_beta_r_backscat:dpl_py_binding = "profiles.inv.atten_beta_a_backscat" ;
	float profile_circular_depol(profile_time,altitude) ;
		profile_circular_depol:long_name = "Circular depolarization ratio profile for particulate" ;
		profile_circular_depol:description = "left circular return divided by right circular return" ;
		profile_circular_depol:units = " " ;
		profile_circular_depol:missing_value = 9.96920996838687e+36 ;
		profile_circular_depol:plot_scale = "logarithmic" ;
		profile_circular_depol:dpl_py_binding = "profiles.inv.circular_depol" ;
	float profile_linear_depol(profile_time,altitude) ;
		profile_linear_depol:long_name = "Linear depolarization ratio profile for particulate" ;
		profile_linear_depol:description = "??? return" ;
		profile_linear_depol:units = " " ;
		profile_linear_depol:missing_value = 9.96920996838687e+36 ;
		profile_linear_depol:plot_scale = "logarithmic" ;
		profile_linear_depol:dpl_py_binding = "profiles.inv.linear_depol" ;
	float profile_molecular_counts(profile_time,altitude) ;
		profile_molecular_counts:long_name = "Molecular Photon Counts profile" ;
		profile_molecular_counts:description = "Raw counts, per averaging interval with pileup, afterpulse, and darkcount corrections applied" ;
		profile_molecular_counts:units = "counts" ;
		profile_molecular_counts:missing_value = -1 ;
		profile_molecular_counts:plot_scale = "logarithmic" ;
		profile_molecular_counts:dpl_py_binding = "profiles.molecular_counts" ;
	float profile_molecular_i2a_counts(profile_time,altitude) ;
		profile_molecular_i2a_counts:long_name = "Molecular I2A Photon Counts profile" ;
		profile_molecular_i2a_counts:description = "Raw counts, per averaging interval with pileup, afterpulse, and darkcount corrections applied" ;
		profile_molecular_i2a_counts:units = "counts" ;
		profile_molecular_i2a_counts:missing_value = -1 ;
		profile_molecular_i2a_counts:plot_scale = "logarithmic" ;
		profile_molecular_i2a_counts:dpl_py_binding = "profiles.molecular_i2a_counts" ;
	float profile_combined_counts_lo(profile_time,altitude) ;
		profile_combined_counts_lo:long_name = "Low Gain Combined Photon Counts profile" ;
		profile_combined_counts_lo:description = "Raw counts, per averaging interval with pileup, afterpulse, and darkcount corrections applied" ;
		profile_combined_counts_lo:units = "counts" ;
		profile_combined_counts_lo:missing_value = -1 ;
		profile_combined_counts_lo:plot_scale = "logarithmic" ;
		profile_combined_counts_lo:dpl_py_binding = "profiles.combined_lo_counts" ;
	float profile_combined_counts_hi(profile_time,altitude) ;
		profile_combined_counts_hi:long_name = "High Gain Combined Photon Counts profile" ;
		profile_combined_counts_hi:description = "Raw counts, per averaging interval with pileup, afterpulse, and darkcount corrections applied" ;
		profile_combined_counts_hi:units = "counts" ;
		profile_combined_counts_hi:missing_value = -1 ;
		profile_combined_counts_hi:plot_scale = "logarithmic" ;
		profile_combined_counts_hi:dpl_py_binding = "profiles.combined_hi_counts" ;
	float profile_cross_counts(profile_time,altitude) ;
		profile_cross_counts:long_name = "Cross Polarized Photon Counts profile" ;
		profile_cross_counts:description = "Raw counts, per averaging interval with pileup, afterpulse, and darkcount corrections applied" ;
		profile_cross_counts:units = "counts" ;
		profile_cross_counts:missing_value = -1 ;
		profile_cross_counts:plot_scale = "logarithmic" ;
		profile_cross_counts:dpl_py_binding = "profiles.cross_pol_counts" ;
	float profile_beta_a_backscat_parallel(profile_time,altitude) ;
		profile_beta_a_backscat_parallel:long_name = "Particulate nondepolarized backscatter cross section profile" ;
		profile_beta_a_backscat_parallel:units = "1/(m sr)" ;
		profile_beta_a_backscat_parallel:missing_value = 9.96920996838687e+36 ;
		profile_beta_a_backscat_parallel:plot_scale = "logarithmic" ;
		profile_beta_a_backscat_parallel:dpl_py_binding = "profiles.inv.beta_a_backscat_par" ;
	float profile_beta_a_backscat(profile_time,altitude) ;
		profile_beta_a_backscat:long_name = "Particulate backscatter cross section profile" ;
		profile_beta_a_backscat:units = "1/(m sr)" ;
		profile_beta_a_backscat:missing_value = 9.96920996838687e+36 ;
		profile_beta_a_backscat:plot_scale = "logarithmic" ;
		profile_beta_a_backscat:dpl_py_binding = "profiles.inv.beta_a_backscat" ;
	float profile_beta_m(altitude) ;
		profile_beta_m:long_name = "Raob molecular scattering cross section profile" ;
		profile_beta_m:units = "1/meter" ;
		profile_beta_m:plot_scale = "logarithmic" ;
		profile_beta_m:dpl_py_binding = "rs_inv.beta_r_backscat" ;
	float profile_Na(profile_time,altitude) ;
		profile_Na:long_name = "Inverted Aerosol Profile" ;
		profile_Na:units = " " ;
		profile_Na:dpl_py_binding = "profiles.inv.Na" ;
	float profile_Nm(profile_time,altitude) ;
		profile_Nm:long_name = "Inverted Molecular Profile" ;
		profile_Nm:units = " " ;
		profile_Nm:dpl_py_binding = "profiles.inv.Nm" ;
	float profile_Nm_i2a(profile_time,altitude) ;
		profile_Nm_i2a:long_name = "Inverted I2A Molecular Profile" ;
		profile_Nm_i2a:units = " " ;
		profile_Nm_i2a:dpl_py_binding = "profiles.inv.Nm_i2a" ;
	float profile_Ncp(profile_time,altitude) ;
		profile_Ncp:long_name = "Inverted Cross Polarization Profile" ;
		profile_Ncp:units = " " ;
		profile_Ncp:dpl_py_binding = "profiles.inv.Ncp" ;

// global attributes:
                :dpl_py_template = "segment_hsrl_profiles.cdl" ;
                :dpl_py_template_version = 20140216 ;
		:time_zone = "UTC" ;
}
