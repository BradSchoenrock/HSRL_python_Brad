netcdf out {
dimensions:
	time = UNLIMITED ;
	altitude = 0 ;
	bin_range = 0 ;
    profile_time = 1;
	time_vector = 8 ;
	calibration = UNLIMITED ; 
	githash = 40;
	sondenamelength = 32 ;
	i2header = 2000 ;
	geoheader = 2000 ;
	apheader = 2000 ;
variables:
	int base_time ;
		base_time:string = "2006-10-23 18:19:59 UTC" ;
		base_time:long_name = "Base seconds since Unix Epoch" ;
		base_time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		base_time:dpl_py_binding = "dne" ;
	short first_time(time_vector) ;
		first_time:long_name = "First Time in file" ;
		first_time:dpl_py_binding = "dne" ;
	short last_time(time_vector) ;
		last_time:long_name = "Last Time in file" ;
		last_time:dpl_py_binding = "dne" ;
	double time(time) ;
		time:long_name = "Time" ;
		time:units = "seconds since 2006-10-23 18:19:59 UTC" ;
		time:dpl_py_binding = "rs_inv.times" ;
        time:dpl_py_type = "python_datetime" ;
	float latitude(time) ;
		latitude:long_name = "latitude of lidar" ;
		latitude:units = "degree_N" ;
		latitude:dpl_py_binding = "rs_mean.latitude" ;
	float longitude(time) ;
		longitude:long_name = "longitude of lidar" ;
		longitude:units = "degree_E" ;
		longitude:dpl_py_binding = "rs_mean.longitude" ;
	float lidar_altitude(time) ;
		lidar_altitude:long_name = "ground based platform altitude" ;
		lidar_altitude:units = "meters" ;
		lidar_altitude:dpl_py_binding = "rs_mean.GPS_MSL_Alt" ;
    float telescope_roll_angle_offset(time) ;
		telescope_roll_angle_offset:long_name = "Telescope Mounting Roll Angle Offset" ;
		telescope_roll_angle_offset:description = "Telescope Mount Roll Angle Relative to platform or aircraft measured clockwise from up" ;
		telescope_roll_angle_offset:units = "degrees" ;
		telescope_roll_angle_offset:range = -180.0, 360.0 ;
		telescope_roll_angle_offset:dpl_py_binding = "rs_mean.telescope_roll_angle_offset" ;
	double sonde_times(calibration) ;
		sonde_times:long_name = "Time of Temperature Profiles" ;
		sonde_times:description = "New raob data" ;
		sonde_times:dpl_py_binding = "sounding.times" ;
        sonde_times:dpl_py_type = "python_datetime" ;
	double sonde_longitude(calibration) ;
		sonde_longitude:long_name = "Longitude of Temperature Profiles" ;
		sonde_longitude:units = "degree_E" ;
		sonde_longitude:description = "Sounding Longitude source" ;
		sonde_longitude:dpl_py_binding = "sounding.longitude" ;
	double sonde_latitude(calibration) ;
		sonde_latitude:long_name = "Latituide of Temperature Profiles" ;
		sonde_latitude:units = "degree_N" ;
		sonde_latitude:description = "Sounding Latitude source" ;
		sonde_latitude:dpl_py_binding = "sounding.latitude" ;
	double new_cal_times(calibration) ;
		new_cal_times:long_name = "Time of Calibration Change" ;
		new_cal_times:description = "New raob or system calibration data triggered recalibration" ;
		new_cal_times:dpl_py_binding = "chunk_start_time" ;
        new_cal_times:dpl_py_type = "python_datetime" ;
	float altitude(altitude) ;
		altitude:long_name = "Height above lidar" ;
		altitude:units = "meters" ;
		altitude:dpl_py_binding = "rs_mean.msl_altitudes" ;
	byte new_cal_trigger(calibration) ;
		new_cal_trigger:long_name = "Trigger of Calibration Change" ;
		new_cal_trigger:description = "reason for recalibration" ;
		new_cal_trigger:bit_0 = "radiosonde profile" ;
		new_cal_trigger:bit_1 = "i2 scan" ;
		new_cal_trigger:bit_2 = "geometry" ;
		new_cal_trigger:dpl_py_required = 1 ;
	short new_cal_offset(calibration) ;
		new_cal_offset:long_name = "Record Dimension equivalent Offset" ;
		new_cal_offset:min_value = 0 ;
		new_cal_offset:dpl_py_binding = "dne" ;
	float top_alt_sounding(calibration) ;
		top_alt_sounding:long_name = "Sounding Maximum Altitude" ;
		top_alt_sounding:units = "meters" ;
		top_alt_sounding:dpl_py_binding = "sounding.top" ;
	float temperature_profile(calibration, altitude) ;
		temperature_profile:long_name = "Raob Temperature Profile" ;
		temperature_profile:description = "Temperature interpolated to requested altitude resolution" ;
		temperature_profile:units = "degrees Kelvin" ;
		temperature_profile:dpl_py_binding = "sounding.temps" ;
	float pressure_profile(calibration,altitude) ;
		pressure_profile:long_name = "Raob pressure Profile" ;
		pressure_profile:description = "Pressure interpolated to requested altitude resolution" ;
		pressure_profile:units = "hectopascals" ;
		pressure_profile:dpl_py_binding = "sounding.pressures" ;
	float dewpoint_profile(calibration, altitude) ;
		dewpoint_profile:long_name = "Raob Dewpoint Temperature Profile" ;
		dewpoint_profile:description = "Dewpoint interpolated to requested altitude resolution" ;
		dewpoint_profile:units = "degrees Kelvin" ;
		dewpoint_profile:missing_value = NaNf ;
		dewpoint_profile:dpl_py_binding = "sounding.dew_points" ;
	float windspeed_profile(calibration, altitude) ;
		windspeed_profile:long_name = "Raob Wind Speed Profile" ;
		windspeed_profile:description = "Speeds interpolated to requested altitude resolution" ;
		windspeed_profile:units = "m/s" ;
		windspeed_profile:missing_value = NaNf ;
		windspeed_profile:dpl_py_binding = "sounding.wind_spd" ;
	float winddir_profile(calibration, altitude) ;
		winddir_profile:long_name = "Raob Wind Direction Profile" ;
		winddir_profile:description = "Directions interpolated to requested altitude resolution" ;
		winddir_profile:units = "degrees" ;
		winddir_profile:missing_value = NaNf ;
		winddir_profile:dpl_py_binding = "sounding.wind_dir" ;
	char calibration_version(calibration, githash) ;
		calibration_version:long_name = "Calibration Tables GIT Version" ;
		calibration_version:dpl_py_binding = "gitversion" ;
	short raob_time_vector(calibration,time_vector) ;
		raob_time_vector:dpl_py_require = 1 ;
	float range_resolution ;
		range_resolution:dpl_py_require = 1 ;
	float time_average ;
		time_average:dpl_py_require = 1 ;
	char raob_station(calibration, sondenamelength) ;
		raob_station:long_name = "Radiosonde Station ID" ;
		raob_station:dpl_py_binding = "sounding.sounding_id" ;
	char i2_txt_header(calibration, i2header) ;
		i2_txt_header:long_name = "i2_scan_file_text_info" ;
		i2_txt_header:description = "Contains name of file used to compute calibration" ;
		i2_txt_header:dpl_py_binding = "rs_cal.i2scan.header" ;
	char geo_txt_header(calibration, geoheader) ;
		geo_txt_header:long_name = "geometric_correction_file_txt_header." ;
		geo_txt_header:dpl_py_binding = "rs_cal.geo.header" ;
	char ap_txt_header(calibration, apheader) ;
		ap_txt_header:long_name = "afterpulse_correction_file_txt_header." ;
		ap_txt_header:dpl_py_binding = "rs_cal.afterpulse.header" ;
	float Cmc(calibration, altitude) ;
		Cmc:long_name = "Molecular in Combined Calibration" ;
		Cmc:dpl_py_binding = "rs_Cxx.Cmc" ;
	float Cmm(calibration, altitude) ;
		Cmm:long_name = "Molecular in Molecular Calibration" ;
		Cmm:dpl_py_binding = "rs_Cxx.Cmm" ;
	float Cam(calibration) ;
		Cam:long_name = "Aerosol in Molecular Calibration" ;
		Cam:dpl_py_binding = "rs_Cxx.Cam" ;
	float Cmm_i2a(calibration, altitude) ;
		Cmm_i2a:long_name = "Molecular in Molecular Calibration" ;
		Cmm_i2a:dpl_py_binding = "rs_Cxx.Cmm_i2a" ;
	float beta_m(calibration, altitude) ;
		beta_m:long_name = "Raob molecular scattering cross section per unit volume" ;
		beta_m:units = "1/meter" ;
		beta_m:plot_scale = "logarithmic" ;
		beta_m:dpl_py_binding = "rs_Cxx.beta_r" ;
	float transmitted_energy(time) ;
		transmitted_energy:long_name = "Transmitted Energy" ;
		transmitted_energy:units = "Joules" ;
		transmitted_energy:missing_value = NaNf ;
		transmitted_energy:dpl_py_binding = "rs_mean.transmitted_energy" ;
	float piezovoltage(time) ;
		piezovoltage:long_name = "piezovoltage" ;
		piezovoltage:units = "Volts" ;
		piezovoltage:missing_value = NaNf ;
		piezovoltage:dpl_py_require = 1 ;
	int num_seeded_shots(time) ;
		num_seeded_shots:long_name = "Number of Seeded Shots" ;
		num_seeded_shots:missing_value = -1 ;
		num_seeded_shots:dpl_py_binding = "rs_mean.seeded_shots" ;
	int num_shots(time) ;
		num_shots:long_name = "Number of Shots" ;
		num_shots:missing_value = -1 ;
		num_shots:dpl_py_binding = "rs_mean.shot_count" ;
	float seed_quality(time) ;
		seed_quality:long_name = "Laser Seeding Quality" ;
		seed_quality:description = "The ratio of seeded shots to total shots. Only seeded shot data is stored and processed.  A low seed ratio can result in low noise resistance." ;
		seed_quality:missing_value = NaNf ;
		seed_quality:range = 0., 1. ;
		seed_quality:dpl_py_require = 1 ;
	float frequency_quality(time) ;
		frequency_quality:long_name = "Laser Frequency Quality" ;
		frequency_quality:description = "An ratio average of how good the frequency lock is per raw interval. A low value can result in poor separation of molecular and aerosol counts." ;
		frequency_quality:missing_value = NaNf ;
		frequency_quality:range = 0., 1. ;
		frequency_quality:dpl_py_require = 1 ;
	float lock_quality(time) ;
		lock_quality:long_name = "Laser Lock Quality" ;
		lock_quality:description = "A ratio of likely locked intervals (frequency_quality>=.5) to seeded intervals.  A low value can result in poor separation of molecular and aerosol counts." ;
		lock_quality:missing_value = NaNf ;
		lock_quality:range = 0., 1. ;
		lock_quality:dpl_py_require = 1 ;
	float mol_cal_pulse(time) ;
		mol_cal_pulse:long_name = "Molecular calibration pulse" ;
		mol_cal_pulse:description = "Sum of photon counts in the molecular channel due to light scattered with the telescope." ;
		mol_cal_pulse:units = "counts" ;
		mol_cal_pulse:missing_value = NaNf ;
		mol_cal_pulse:dpl_py_binding = "rs_mean.molecular_cal_pulse" ;
	float mol_i2a_cal_pulse(time) ;
		mol_i2a_cal_pulse:long_name = "Molecular I2A calibration pulse" ;
		mol_i2a_cal_pulse:description = "Sum of photon counts in the molecular channel due to light scattered with the telescope." ;
		mol_i2a_cal_pulse:units = "counts" ;
		mol_i2a_cal_pulse:missing_value = NaNf ;
		mol_i2a_cal_pulse:dpl_py_binding = "rs_mean.molecular_i2a_cal_pulse" ;
	int mol_norm_idx ;
		mol_norm_idx:dpl_py_binding = "rs_inv.mol_norm_index" ;
	float c_pol_dark_count(time) ;
		c_pol_dark_count:long_name = "Cross Polarization Dark Count FIXME dark counts need alt" ;
		c_pol_dark_count:description = "Counts/bin at output resolution" ;
		c_pol_dark_count:units = "counts" ;
		c_pol_dark_count:missing_value = NaNf ;
		c_pol_dark_count:dpl_py_binding = "rs_mean.c_pol_dark_counts" ;
	float mol_i2a_dark_count(time) ;
		mol_i2a_dark_count:long_name = "Molecular I2A Dark Count" ;
		mol_i2a_dark_count:description = "Counts/bin at output resolution" ;
		mol_i2a_dark_count:units = "counts" ;
		mol_i2a_dark_count:missing_value = NaNf ;
		mol_i2a_dark_count:dpl_py_binding = "rs_mean.mol_i2a_dark_counts" ;
	float mol_dark_count(time) ;
		mol_dark_count:long_name = "Molecular Dark Count" ;
		mol_dark_count:description = "Counts/bin at output resolution" ;
		mol_dark_count:units = "counts" ;
		mol_dark_count:missing_value = NaNf ;
		mol_dark_count:dpl_py_binding = "rs_mean.mol_dark_counts" ;
	float combined_dark_count_lo(time) ;
		combined_dark_count_lo:long_name = "Low Gain Combined Dark Count" ;
		combined_dark_count_lo:description = "Counts/bin at output resolution" ;
		combined_dark_count_lo:units = "counts" ;
		combined_dark_count_lo:missing_value = NaNf ;
		combined_dark_count_lo:dpl_py_binding = "rs_mean.c_lo_dark_counts" ;
	float combined_dark_count_hi(time) ;
		combined_dark_count_hi:long_name = "High Gain Combined Dark Count" ;
		combined_dark_count_hi:description = "Counts/bin at output resolution" ;
		combined_dark_count_hi:units = "counts" ;
		combined_dark_count_hi:missing_value = NaNf ;
		combined_dark_count_hi:dpl_py_binding = "rs_mean.c_hi_dark_counts" ;
	float combined_1064_dark_count(time) ;
		combined_1064_dark_count:long_name = "Combined 1064 Dark Count" ;
		combined_1064_dark_count:description = "Counts/bin at output resolution" ;
		combined_1064_dark_count:units = "counts" ;
		combined_1064_dark_count:missing_value = NaNf ;
		combined_1064_dark_count:dpl_py_binding = "rs_mean.combined_1064_dark_count" ;
	float combined_dark_count(time) ;
		combined_dark_count:long_name = "Combined Dark Count" ;
		combined_dark_count:description = "Counts/bin at output resolution" ;
		combined_dark_count:units = "counts" ;
		combined_dark_count:missing_value = NaNf ;
		combined_dark_count:dpl_py_binding = "rs_mean.c_dark_counts" ;
	float combined_gain(calibration) ;
		combined_gain:long_name = "Combined Gain Factor" ;
		combined_gain:description = "Low Gain level * Factor ~ High Gain level" ;
		combined_gain:dpl_py_binding = "rs_constants.hi_to_low_combined_channel_gain_ratio" ;
	float combined_merge_threshhold(calibration) ;
		combined_merge_threshhold:long_name = "Combined Merge Threshhold" ;
		combined_merge_threshhold:dpl_py_binding = "rs_constants.combined_channel_merge_threshhold" ;
	float polarization_cross_talk(calibration) ;
		polarization_cross_talk:long_name = "Polarization Cross Talk" ;
		polarization_cross_talk:dpl_py_binding = "rs_constants.polarization_cross_talk" ;
	float wfov_to_combined_gain_ratio(calibration) ;
		wfov_to_combined_gain_ratio:long_name = "WFOV to Combined Gain" ;
		wfov_to_combined_gain_ratio:dpl_py_binding = "rs_constants.wfov_to_combined_gain_ratio" ;
	float combined_to_cross_pol_gain_ratio(calibration) ;
		combined_to_cross_pol_gain_ratio:long_name = "Combined to Cross Pol Gain" ;
		combined_to_cross_pol_gain_ratio:dpl_py_binding = "rs_constants.combined_to_cross_pol_gain_ratio" ;
	float molecular_to_wfov_gain_ratio(calibration) ;
		molecular_to_wfov_gain_ratio:long_name = "Molecular to WFOV Gain" ;
		molecular_to_wfov_gain_ratio:dpl_py_binding = "rs_constants.molecular_to_wfov_gain_ratio" ;
	float geo_cor(calibration, bin_range) ;
		geo_cor:long_name = "Overlap correction" ;
		geo_cor:description = "Geometric overlap correction in raw range bins" ;
		geo_cor:units = " " ;
		geo_cor:missing_value = NaNf ;
		geo_cor:plot_scale = "logarithmic" ;
		geo_cor:dpl_py_binding = "geo_corr" ;
	int od_norm_index ;
		od_norm_index:long_name = "Optical depth normalization index FIXME shouldn't be needed" ;
		od_norm_index:description = "optical depth reference bin. normalized so Optical Depth is 0 at this altitude index" ;
		od_norm_index:dpl_py_binding = "rs_inv.od_norm_index" ;
	float od(time, altitude) ;
		od:long_name = "Aerosol + Molecular Optical Depth" ;
		od:units = " " ;
		od:missing_value = NaNf ;
		od:insufficient_data = NaNf ;
		od:plot_scale = "logarithmic" ;
		od:dpl_py_binding = "rs_inv.optical_depth" ;
	float profile_temperature(profile_time,altitude) ;
		profile_temperature:long_name = "HSRL I2A Temperature Profile" ;
		profile_temperature:description = "HSRL Temperature Profile derived the comparison of I2A to I2 filtered molecular channels" ;
		profile_temperature:units = "degK" ;
		profile_temperature:missing_value = NaNf ;
		profile_temperature:insufficient_data = NaNf ;
		profile_temperature:dpl_py_binding = "profiles.i2a_temperatures" ;
	float profile_od(profile_time,altitude) ;
		profile_od:long_name = "Aerosol + Molecular Optical Depth Profile" ;
		profile_od:units = " " ;
		profile_od:missing_value = NaNf ;
		profile_od:insufficient_data = NaNf ;
		profile_od:plot_scale = "logarithmic" ;
		profile_od:dpl_py_binding = "profiles.inv.optical_depth" ;
	float profile_extinction(profile_time,altitude) ;
		profile_extinction:long_name = "Aerosol + Molecular Extinction Profile" ;
		profile_extinction:units = " " ;
		profile_extinction:missing_value = NaNf ;
		profile_extinction:insufficient_data = NaNf ;
		profile_extinction:plot_scale = "logarithmic" ;
		profile_extinction:dpl_py_binding = "profiles.inv.extinction" ;
	float extinction(time,altitude) ;
		extinction:long_name = "Aerosol + Molecular Extinction Profile" ;
		extinction:units = " " ;
		extinction:missing_value = NaNf ;
		extinction:insufficient_data = NaNf ;
		extinction:plot_scale = "logarithmic" ;
		extinction:dpl_py_binding = "rs_inv.extinction" ;
	float od_aerosol(time, altitude) ;
		od_aerosol:long_name = "Aerosol Optical Depth" ;
		od_aerosol:units = " " ;
		od_aerosol:missing_value = NaNf ;
		od_aerosol:insufficient_data = NaNf ;
		od_aerosol:plot_scale = "logarithmic" ;
		od_aerosol:dpl_py_binding = "rs_inv.optical_depth_aerosol" ;
	float profile_od_aerosol(profile_time,altitude) ;
		profile_od_aerosol:long_name = "Aerosol Optical Depth Profile" ;
		profile_od_aerosol:units = " " ;
		profile_od_aerosol:missing_value = NaNf ;
		profile_od_aerosol:insufficient_data = NaNf ;
		profile_od_aerosol:plot_scale = "logarithmic" ;
		profile_od_aerosol:dpl_py_binding = "profiles.inv.optical_depth_aerosol" ;
	float profile_extinction_aerosol(profile_time,altitude) ;
		profile_extinction_aerosol:long_name = "Aerosol Extinction Profile" ;
		profile_extinction_aerosol:units = " " ;
		profile_extinction_aerosol:missing_value = NaNf ;
		profile_extinction_aerosol:insufficient_data = NaNf ;
		profile_extinction_aerosol:plot_scale = "logarithmic" ;
		profile_extinction_aerosol:dpl_py_binding = "profiles.inv.extinction_aerosol" ;
	float extinction_aerosol(time,altitude) ;
		extinction_aerosol:long_name = "Aerosol Extinction" ;
		extinction_aerosol:units = " " ;
		extinction_aerosol:missing_value = NaNf ;
		extinction_aerosol:insufficient_data = NaNf ;
		extinction_aerosol:plot_scale = "logarithmic" ;
		extinction_aerosol:dpl_py_binding = "rs_inv.extinction_aerosol" ;
	float radar_backscattercrosssection(time, altitude) ;
		radar_backscattercrosssection:long_name = "Radar Backscatter Cross Section" ;
		radar_backscattercrosssection:units = "1/(m sr)" ;
		radar_backscattercrosssection:missing_value = NaNf ;
		radar_backscattercrosssection:dpl_py_binding = "rs_mmcr.Backscatter" ;
	float radar_reflectivity(time, altitude) ;
		radar_reflectivity:long_name = "Radar Reflectivity" ;
		radar_reflectivity:units = "dBz" ;
		radar_reflectivity:missing_value = NaNf ;
		radar_reflectivity:dpl_py_binding = "rs_mmcr.Reflectivity" ;
	float radar_spectralwidth(time, altitude) ;
		radar_spectralwidth:long_name = "Radar Spectral Width" ;
		radar_spectralwidth:units = "m/s" ;
		radar_spectralwidth:missing_value = NaNf ;
		radar_spectralwidth:dpl_py_binding = "rs_mmcr.SpectralWidth" ;
	float radar_dopplervelocity(time, altitude) ;
		radar_dopplervelocity:long_name = "Radar doppler Velocity" ;
		radar_dopplervelocity:units = "m/s" ;
		radar_dopplervelocity:missing_value = NaNf ;
		radar_dopplervelocity:dpl_py_binding = "rs_mmcr.MeanDopplerVelocity" ;
	float effective_diameter_prime(time, altitude) ;
		effective_diameter_prime:long_name = "lidar/radar effective particle diameter prime measurement" ;
		effective_diameter_prime:units = "m" ;
		effective_diameter_prime:description = "Effective diameter directly from the ratio of Lidar Backscatter and Radar Reflectivity; (<volume^2>/<area>)^.25, see Donovan JGR Nov 2001" ;
		effective_diameter_prime:missing_value = NaNf ;
		effective_diameter_prime:dpl_py_binding = "rs_spheroid_particle.effective_diameter_prime" ;
	float effective_diameter(time, altitude) ;
		effective_diameter:long_name = "Effective particle diameter" ;
		effective_diameter:units = "m" ;
		effective_diameter:description = "Effective particle diameter derived from ratio of Lidar Backscatter and Radar Reflectivity; assuming a gamma size distribution using assumptions from particle processing parameters" ;
		effective_diameter:missing_value = NaNf ;
		effective_diameter:dpl_py_binding = "rs_spheroid_particle.effective_diameter" ;
	float num_particles(time, altitude) ;
		num_particles:long_name = "Number density of particles" ;
		num_particles:units = "1/liter" ;
		num_particles:description = "Number of particles per liter derived from ratio of lidar backscatter and radar reflectivity; assuming a gamma size distribution" ;
		num_particles:missing_value = NaNf ;
		num_particles:dpl_py_binding = "rs_spheroid_particle.num_particles" ;
	float mean_diameter(time, altitude) ;
		mean_diameter:long_name = "Mean diameter of particles" ;
		mean_diameter:units = "m" ;
		mean_diameter:description = "Mean diameter of particles derived from the effective diameter and the gamma size distribution" ;
		mean_diameter:missing_value = NaNf ;
		mean_diameter:dpl_py_binding = "rs_spheroid_particle.mean_diameter" ;
	float LWC(time, altitude) ;
		LWC:long_name = "Liquid water content" ;
		LWC:units = "kg/m^3" ;
		LWC:description = "Liquid water content derived from ratio of lidar backscatter and radar reflectivity; assuming a gamma size distribution" ;
		LWC:missing_value = NaNf ;
		LWC:dpl_py_binding = "rs_spheroid_particle.LWC" ;
	float precip_rate(time, altitude) ;
		precip_rate:long_name = "HSRL-Radar Precipitation Rate" ;
		precip_rate:units = "m/s" ;
		precip_rate:description = "precipitation accumulation rate from combined hsrl radar retrieval" ;
		precip_rate:missing_value = NaNf ;
		precip_rate:dpl_py_binding = "rs_spheroid_particle.hsrl_radar_precip_rate" ;
	float fall_velocity(time, altitude) ;
		fall_velocity:long_name = "radar-weighted fall velocity" ;
		fall_velocity:units = "m/s" ;
		fall_velocity:description = "modeled fall velocity weighted by radar cross section" ;
		fall_velocity:missing_value = NaNf ;
		fall_velocity:dpl_py_binding = "rs_spheroid_particle.rw_fall_velocity" ;
	float model_spectral_width(time, altitude) ;
		model_spectral_width:long_name = "Modeled Radar Spectral Width" ;
		model_spectral_width:units = "m/s" ;
		model_spectral_width:description = "radar spectral width modeled from derived hsrl_radar particle size retrieval" ;
		model_spectral_width:missing_value = NaNf ;
		model_spectral_width:dpl_py_binding = "rs_spheroid_particle.model_spectral_width" ;
	float atten_beta_r_backscat(time, altitude) ;
		atten_beta_r_backscat:long_name = "Attenuated Molecular return" ;
		atten_beta_r_backscat:units = "1/(m sr)" ;
		atten_beta_r_backscat:missing_value = NaNf ;
		atten_beta_r_backscat:plot_scale = "logarithmic" ;
		atten_beta_r_backscat:dpl_py_binding = "rs_inv.atten_beta_a_backscat" ;
	float profile_atten_beta_r_backscat(altitude) ;
		profile_atten_beta_r_backscat:long_name = "Attenuated Molecular Profile" ;
		profile_atten_beta_r_backscat:units = "1/(m sr)" ;
		profile_atten_beta_r_backscat:missing_value = NaNf ;
		profile_atten_beta_r_backscat:plot_scale = "logarithmic" ;
		profile_atten_beta_r_backscat:dpl_py_binding = "profiles.inv.atten_beta_a_backscat" ;
	float circular_depol(time, altitude) ;
		circular_depol:long_name = "Circular depolarization ratio for particulate" ;
		circular_depol:description = "left circular return divided by right circular return" ;
		circular_depol:units = " " ;
		circular_depol:missing_value = NaNf ;
		circular_depol:plot_scale = "logarithmic" ;
		circular_depol:dpl_py_binding = "rs_inv.circular_depol" ;
	float linear_depol(time, altitude) ;
		linear_depol:long_name = "Linear depolarization ratio for particulate" ;
		linear_depol:description = "Perpendicular / parallel polarization" ;
		linear_depol:units = " " ;
		linear_depol:missing_value = NaNf ;
		linear_depol:plot_scale = "logarithmic" ;
		linear_depol:dpl_py_binding = "rs_inv.linear_depol" ;
	float profile_circular_depol(profile_time,altitude) ;
		profile_circular_depol:long_name = "Circular depolarization ratio profile for particulate" ;
		profile_circular_depol:description = "left circular return divided by right circular return" ;
		profile_circular_depol:units = " " ;
		profile_circular_depol:missing_value = NaNf ;
		profile_circular_depol:plot_scale = "logarithmic" ;
		profile_circular_depol:dpl_py_binding = "profiles.inv.circular_depol" ;
	float profile_linear_depol(profile_time,altitude) ;
		profile_linear_depol:long_name = "Linear depolarization ratio profile for particulate" ;
		profile_linear_depol:description = "Perpendicular / parallel polarization" ;
		profile_linear_depol:units = " " ;
		profile_linear_depol:missing_value = NaNf ;
		profile_linear_depol:plot_scale = "logarithmic" ;
		profile_linear_depol:dpl_py_binding = "profiles.inv.linear_depol" ;
	float profile_molecular_counts(profile_time,altitude) ;
		profile_molecular_counts:long_name = "Molecular Photon Counts profile" ;
		profile_molecular_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		profile_molecular_counts:units = "counts" ;
		profile_molecular_counts:missing_value = NaNf ;
		profile_molecular_counts:plot_scale = "logarithmic" ;
		profile_molecular_counts:dpl_py_binding = "profiles.molecular_counts" ;
	float profile_molecular_i2a_counts(profile_time,altitude) ;
		profile_molecular_i2a_counts:long_name = "Molecular I2A Photon Counts profile" ;
		profile_molecular_i2a_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		profile_molecular_i2a_counts:units = "counts" ;
		profile_molecular_i2a_counts:missing_value = NaNf ;
		profile_molecular_i2a_counts:plot_scale = "logarithmic" ;
		profile_molecular_i2a_counts:dpl_py_binding = "profiles.molecular_i2a_counts" ;
	float profile_combined_counts_lo(profile_time,altitude) ;
		profile_combined_counts_lo:long_name = "Low Gain Combined Photon Counts profile" ;
		profile_combined_counts_lo:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		profile_combined_counts_lo:units = "counts" ;
		profile_combined_counts_lo:missing_value = NaNf ;
		profile_combined_counts_lo:plot_scale = "logarithmic" ;
		profile_combined_counts_lo:dpl_py_binding = "profiles.combined_lo_counts" ;
	float profile_combined_counts_hi(profile_time,altitude) ;
		profile_combined_counts_hi:long_name = "High Gain Combined Photon Counts profile" ;
		profile_combined_counts_hi:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		profile_combined_counts_hi:units = "counts" ;
		profile_combined_counts_hi:missing_value = NaNf ;
		profile_combined_counts_hi:plot_scale = "logarithmic" ;
		profile_combined_counts_hi:dpl_py_binding = "profiles.combined_hi_counts" ;
	float profile_combined_counts(profile_time,altitude) ;
		profile_combined_counts:long_name = "Combined Photon Counts profile" ;
		profile_combined_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		profile_combined_counts:units = "counts" ;
		profile_combined_counts:missing_value = NaNf ;
		profile_combined_counts:plot_scale = "logarithmic" ;
		profile_combined_counts:dpl_py_binding = "profiles.combined_counts" ;
	float profile_combined_1064_counts(profile_time,altitude) ;
		profile_combined_1064_counts:long_name = "Combined 1064nm Photon Counts profile" ;
		profile_combined_1064_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		profile_combined_1064_counts:units = "counts" ;
		profile_combined_1064_counts:missing_value = NaNf ;
		profile_combined_1064_counts:plot_scale = "logarithmic" ;
		profile_combined_1064_counts:dpl_py_binding = "profiles.combined_1064_counts" ;
	float profile_cross_counts(profile_time,altitude) ;
		profile_cross_counts:long_name = "Cross Polarized Photon Counts profile" ;
		profile_cross_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		profile_cross_counts:units = "counts" ;
		profile_cross_counts:missing_value = NaNf ;
		profile_cross_counts:plot_scale = "logarithmic" ;
		profile_cross_counts:dpl_py_binding = "profiles.cross_pol_counts" ;
	float profile_molecular_raw_counts(profile_time,altitude) ;
		profile_molecular_raw_counts:long_name = "Molecular Raw Photon Counts profile" ;
		profile_molecular_raw_counts:description = "Raw counts profile with pileup correction applied" ;
		profile_molecular_raw_counts:units = "counts" ;
		profile_molecular_raw_counts:missing_value = NaNf ;
		profile_molecular_raw_counts:plot_scale = "logarithmic" ;
		profile_molecular_raw_counts:dpl_py_binding = "profiles.raw_molecular_counts" ;
	float profile_molecular_i2a_raw_counts(profile_time,altitude) ;
		profile_molecular_i2a_raw_counts:long_name = "Molecular I2A Raw Photon Counts profile" ;
		profile_molecular_i2a_raw_counts:description = "Raw counts profile with pileup correction applied" ;
		profile_molecular_i2a_raw_counts:units = "counts" ;
		profile_molecular_i2a_raw_counts:missing_value = NaNf ;
		profile_molecular_i2a_raw_counts:plot_scale = "logarithmic" ;
		profile_molecular_i2a_raw_counts:dpl_py_binding = "profiles.raw_molecular_i2a_counts" ;
	float profile_combined_raw_counts_lo(profile_time,altitude) ;
		profile_combined_raw_counts_lo:long_name = "Low Gain Combined Raw Photon Counts profile" ;
		profile_combined_raw_counts_lo:description = "Raw counts profile with pileup correction applied" ;
		profile_combined_raw_counts_lo:units = "counts" ;
		profile_combined_raw_counts_lo:missing_value = NaNf ;
		profile_combined_raw_counts_lo:plot_scale = "logarithmic" ;
		profile_combined_raw_counts_lo:dpl_py_binding = "profiles.raw_combined_lo_counts" ;
	float profile_combined_raw_counts_hi(profile_time,altitude) ;
		profile_combined_raw_counts_hi:long_name = "High Gain Combined Raw Photon Counts profile" ;
		profile_combined_raw_counts_hi:description = "Raw counts profile with pileup correction applied" ;
		profile_combined_raw_counts_hi:units = "counts" ;
		profile_combined_raw_counts_hi:missing_value = NaNf ;
		profile_combined_raw_counts_hi:plot_scale = "logarithmic" ;
		profile_combined_raw_counts_hi:dpl_py_binding = "profiles.raw_combined_hi_counts" ;
	float profile_combined_raw_counts(profile_time,altitude) ;
		profile_combined_raw_counts:long_name = "Combined Raw Photon Counts profile" ;
		profile_combined_raw_counts:description = "Raw counts profile with pileup correction applied" ;
		profile_combined_raw_counts:units = "counts" ;
		profile_combined_raw_counts:missing_value = NaNf ;
		profile_combined_raw_counts:plot_scale = "logarithmic" ;
		profile_combined_raw_counts:dpl_py_binding = "profiles.raw_combined_counts" ;
	float profile_combined_wfov_raw_counts(profile_time,altitude) ;
		profile_combined_wfov_raw_counts:long_name = "Combined WFOV Raw Photon Counts profile" ;
		profile_combined_wfov_raw_counts:description = "Raw counts profile with pileup correction applied" ;
		profile_combined_wfov_raw_counts:units = "counts" ;
		profile_combined_wfov_raw_counts:missing_value = NaNf ;
		profile_combined_wfov_raw_counts:plot_scale = "logarithmic" ;
		profile_combined_wfov_raw_counts:dpl_py_binding = "profiles.raw_combined_wfov_counts" ;
	float profile_molecular_wfov_raw_counts(profile_time,altitude) ;
		profile_molecular_wfov_raw_counts:long_name = "Molecular WFOV Raw Photon Counts profile" ;
		profile_molecular_wfov_raw_counts:description = "Raw counts profile with pileup correction applied" ;
		profile_molecular_wfov_raw_counts:units = "counts" ;
		profile_molecular_wfov_raw_counts:missing_value = NaNf ;
		profile_molecular_wfov_raw_counts:plot_scale = "logarithmic" ;
		profile_molecular_wfov_raw_counts:dpl_py_binding = "profiles.raw_molecular_wfov_counts" ;
	float profile_combined_1064_raw_counts(profile_time,altitude) ;
		profile_combined_1064_raw_counts:long_name = "Combined 1064nm Raw Photon Counts profile" ;
		profile_combined_1064_raw_counts:description = "Raw counts profile with pileup correction applied" ;
		profile_combined_1064_raw_counts:units = "counts" ;
		profile_combined_1064_raw_counts:missing_value = NaNf ;
		profile_combined_1064_raw_counts:plot_scale = "logarithmic" ;
		profile_combined_1064_raw_counts:dpl_py_binding = "profiles.raw_combined_1064_counts" ;
	float profile_cross_raw_counts(profile_time,altitude) ;
		profile_cross_raw_counts:long_name = "Cross Polarized Photon Raw Counts profile" ;
		profile_cross_raw_counts:description = "Raw counts profile with pileup correction applied" ;
		profile_cross_raw_counts:units = "counts" ;
		profile_cross_raw_counts:missing_value = NaNf ;
		profile_cross_raw_counts:plot_scale = "logarithmic" ;
		profile_cross_raw_counts:dpl_py_binding = "profiles.raw_cross_pol_counts" ;
	float profile_beta_a_backscat_parallel(profile_time,altitude) ;
		profile_beta_a_backscat_parallel:long_name = "Particulate nondepolarized backscatter cross section profile" ;
		profile_beta_a_backscat_parallel:units = "1/(m sr)" ;
		profile_beta_a_backscat_parallel:missing_value = NaNf ;
		profile_beta_a_backscat_parallel:plot_scale = "logarithmic" ;
		profile_beta_a_backscat_parallel:dpl_py_binding = "profiles.inv.beta_a_backscat_par" ;
	float profile_beta_a_backscat(profile_time,altitude) ;
		profile_beta_a_backscat:long_name = "Particulate backscatter cross section profile" ;
		profile_beta_a_backscat:units = "1/(m sr)" ;
		profile_beta_a_backscat:missing_value = NaNf ;
		profile_beta_a_backscat:plot_scale = "logarithmic" ;
		profile_beta_a_backscat:dpl_py_binding = "profiles.inv.beta_a_backscat" ;
	float beta_a_backscat_parallel(time, altitude) ;
		beta_a_backscat_parallel:long_name = "Particulate nondepolarized backscatter cross section per unit volume" ;
		beta_a_backscat_parallel:units = "1/(m sr)" ;
		beta_a_backscat_parallel:missing_value = NaNf ;
		beta_a_backscat_parallel:plot_scale = "logarithmic" ;
		beta_a_backscat_parallel:dpl_py_binding = "rs_inv.beta_a_backscat_par" ;
	float beta_a(time, altitude) ;
		beta_a:long_name = "Particulate backscatter cross section per unit volume" ;
		beta_a:units = "1/(m sr)" ;
		beta_a:missing_value = NaNf ;
		beta_a:plot_scale = "logarithmic" ;
		beta_a:dpl_py_binding = "rs_inv.beta_a_backscat" ;
	float beta_a_backscat(time, altitude) ;
		beta_a_backscat:long_name = "Particulate backscatter cross section per unit volume" ;
		beta_a_backscat:units = "1/(m sr)" ;
		beta_a_backscat:missing_value = NaNf ;
		beta_a_backscat:plot_scale = "logarithmic" ;
		beta_a_backscat:dpl_py_binding = "rs_inv.beta_a_backscat" ;
	float integrated_backscat(time, altitude) ;
		integrated_backscat:long_name = "Range-integrated backscatter cross section" ;
		integrated_backscat:units = "1/sr" ;
		integrated_backscat:missing_value = NaNf ;
		integrated_backscat:plot_scale = "logarithmic" ;
		integrated_backscat:dpl_py_binding = "rs_inv.integrated_backscatter" ;
	float molecular_counts(time, altitude) ;
		molecular_counts:long_name = "Molecular Photon Counts" ;
		molecular_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		molecular_counts:units = "counts" ;
		molecular_counts:missing_value = NaNf ;
		molecular_counts:plot_scale = "logarithmic" ;
		molecular_counts:dpl_py_binding = "rs_mean.molecular_counts" ;
	float molecular_i2a_counts(time, altitude) ;
		molecular_i2a_counts:long_name = "Molecular I2A Photon Counts" ;
		molecular_i2a_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		molecular_i2a_counts:units = "counts" ;
		molecular_i2a_counts:missing_value = NaNf ;
		molecular_i2a_counts:plot_scale = "logarithmic" ;
		molecular_i2a_counts:dpl_py_binding = "rs_mean.molecular_i2a_counts" ;
	float combined_counts_lo(time, altitude) ;
		combined_counts_lo:long_name = "Low Gain Combined Photon Counts" ;
		combined_counts_lo:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		combined_counts_lo:units = "counts" ;
		combined_counts_lo:missing_value = NaNf ;
		combined_counts_lo:plot_scale = "logarithmic" ;
		combined_counts_lo:dpl_py_binding = "rs_mean.combined_lo_counts" ;
	float combined_counts_hi(time, altitude) ;
		combined_counts_hi:long_name = "High Gain Combined Photon Counts" ;
		combined_counts_hi:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		combined_counts_hi:units = "counts" ;
		combined_counts_hi:missing_value = NaNf ;
		combined_counts_hi:plot_scale = "logarithmic" ;
		combined_counts_hi:dpl_py_binding = "rs_mean.combined_hi_counts" ;
	float combined_1064_counts(time, altitude) ;
		combined_1064_counts:long_name = "Combined 1064nm Photon Counts" ;
		combined_1064_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		combined_1064_counts:units = "counts" ;
		combined_1064_counts:missing_value = NaNf ;
		combined_1064_counts:plot_scale = "logarithmic" ;
		combined_1064_counts:dpl_py_binding = "rs_mean.combined_1064_counts" ;
	float combined_counts(time, altitude) ;
		combined_counts:long_name = "Combined Photon Counts" ;
		combined_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		combined_counts:units = "counts" ;
		combined_counts:missing_value = NaNf ; 
		combined_counts:plot_scale = "logarithmic" ;
		combined_counts:dpl_py_binding = "rs_mean.combined_counts" ;
	float molecular_wfov_counts(time, altitude) ;
		molecular_wfov_counts:long_name = "Molecular WFOV Photon Counts" ;
		molecular_wfov_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		molecular_wfov_counts:units = "counts" ;
		molecular_wfov_counts:missing_value = NaNf ;
		molecular_wfov_counts:plot_scale = "logarithmic" ;
		molecular_wfov_counts:dpl_py_binding = "rs_mean.molecular_wfov_counts" ;
	float combined_wfov_counts(time, altitude) ;
		combined_wfov_counts:long_name = "Combined WFOV Photon Counts" ;
		combined_wfov_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		combined_wfov_counts:units = "counts" ;
		combined_wfov_counts:missing_value = NaNf ;
		combined_wfov_counts:plot_scale = "logarithmic" ;
		combined_wfov_counts:dpl_py_binding = "rs_mean.combined_wfov_counts" ;
	float cross_counts(time, altitude) ;
		cross_counts:long_name = "Cross Polarized Photon Counts" ;
		cross_counts:description = "Raw counts per bin at output resolution with pileup, afterpulse, and darkcount corrections applied" ;
		cross_counts:units = "counts" ;
		cross_counts:missing_value = NaNf ;
		cross_counts:plot_scale = "logarithmic" ;
		cross_counts:dpl_py_binding = "rs_mean.cross_pol_counts" ;
	int molecular_raw_counts(time, altitude) ;
		molecular_raw_counts:long_name = "Molecular Raw Uncorrected Photon Counts" ;
		molecular_raw_counts:description = "Raw counts, per averaging interval with pileup correction applied" ;
		molecular_raw_counts:units = "counts" ;
		molecular_raw_counts:missing_value = -1 ;
		molecular_raw_counts:plot_scale = "logarithmic" ;
		molecular_raw_counts:dpl_py_binding = "rs_mean.raw_molecular_counts" ;
	int molecular_i2a_raw_counts(time, altitude) ;
		molecular_i2a_raw_counts:long_name = "Molecular I2A Raw Uncorrected Photon Counts" ;
		molecular_i2a_raw_counts:description = "Raw counts, per averaging interval with pileup correction applied" ;
		molecular_i2a_raw_counts:units = "counts" ;
		molecular_i2a_raw_counts:missing_value = -1 ;
		molecular_i2a_raw_counts:plot_scale = "logarithmic" ;
		molecular_i2a_raw_counts:dpl_py_binding = "rs_mean.raw_molecular_i2a_counts" ;
	int combined_raw_counts_lo(time, altitude) ;
		combined_raw_counts_lo:long_name = "Low Gain Combined Raw Uncorrected Photon Counts" ;
		combined_raw_counts_lo:description = "Raw counts, per averaging interval with pileup correction applied" ;
		combined_raw_counts_lo:units = "counts" ;
		combined_raw_counts_lo:missing_value = -1 ;
		combined_raw_counts_lo:plot_scale = "logarithmic" ;
		combined_raw_counts_lo:dpl_py_binding = "rs_mean.raw_combined_lo_counts" ;
	int combined_raw_counts_hi(time, altitude) ;
		combined_raw_counts_hi:long_name = "High Gain Combined Raw Uncorrected Photon Counts" ;
		combined_raw_counts_hi:description = "Raw counts, per averaging interval with pileup correction applied" ;
		combined_raw_counts_hi:units = "counts" ;
		combined_raw_counts_hi:missing_value = -1 ;
		combined_raw_counts_hi:plot_scale = "logarithmic" ;
		combined_raw_counts_hi:dpl_py_binding = "rs_mean.raw_combined_hi_counts" ;
	int combined_wfov_raw_counts(time, altitude) ;
		combined_wfov_raw_counts:long_name = "Combined WFOV Raw Uncorrected Photon Counts" ;
		combined_wfov_raw_counts:description = "Raw counts, per averaging interval with pileup correction applied" ;
		combined_wfov_raw_counts:units = "counts" ;
		combined_wfov_raw_counts:missing_value = -1 ;
		combined_wfov_raw_counts:plot_scale = "logarithmic" ;
		combined_wfov_raw_counts:dpl_py_binding = "rs_mean.raw_combined_wfov_counts" ;
	int molecular_wfov_raw_counts(time, altitude) ;
		molecular_wfov_raw_counts:long_name = "Molecular WFOV Raw Uncorrected Photon Counts" ;
		molecular_wfov_raw_counts:description = "Raw counts, per averaging interval with pileup correction applied" ;
		molecular_wfov_raw_counts:units = "counts" ;
		molecular_wfov_raw_counts:missing_value = -1 ;
		molecular_wfov_raw_counts:plot_scale = "logarithmic" ;
		molecular_wfov_raw_counts:dpl_py_binding = "rs_mean.raw_molecular_wfov_counts" ;
	int combined_raw_counts(time, altitude) ;
		combined_raw_counts:long_name = "Combined Raw Uncorrected Photon Counts" ;
		combined_raw_counts:description = "Raw counts, per averaging interval with pileup correction applied" ;
		combined_raw_counts:units = "counts" ;
		combined_raw_counts:missing_value = -1 ;
		combined_raw_counts:plot_scale = "logarithmic" ;
		combined_raw_counts:dpl_py_binding = "rs_mean.raw_combined_counts" ;
	int combined_1064_raw_counts(time, altitude) ;
		combined_1064_raw_counts:long_name = "Combined 1064nm Raw Uncorrected Photon Counts" ;
		combined_1064_raw_counts:description = "Raw counts, per averaging interval with pileup correction applied" ;
		combined_1064_raw_counts:units = "counts" ;
		combined_1064_raw_counts:missing_value = -1 ;
		combined_1064_raw_counts:plot_scale = "logarithmic" ;
		combined_1064_raw_counts:dpl_py_binding = "rs_mean.raw_combined_1064_counts" ;
	int cross_raw_counts(time, altitude) ;
		cross_raw_counts:long_name = "Cross Polarized Raw Uncorrected Photon Counts" ;
		cross_raw_counts:description = "Raw counts, per averaging interval with pileup correction applied" ;
		cross_raw_counts:units = "counts" ;
		cross_raw_counts:missing_value = -1 ;
		cross_raw_counts:plot_scale = "logarithmic" ;
		cross_raw_counts:dpl_py_binding = "rs_mean.raw_cross_pol_counts" ;
	float Na(time, altitude) ;
		Na:long_name = "Range-corrected Number of Aerosol Photons" ;
		Na:description = "Inverted Aerosol times range^2 (in m) divided by 10^6" ;
		Na:units = " " ;
		Na:dpl_py_binding = "rs_inv.Na" ;
	float Nm(time, altitude) ;
		Nm:long_name = "Range-corrected Number of Molecular Photons" ;
		Nm:description = "Inverted Molecular times range^2 (in m) divided by 10^6" ;
		Nm:units = " " ;
		Nm:dpl_py_binding = "rs_inv.Nm" ;
	float Nm_i2a(time, altitude) ;
		Nm_i2a:long_name = "Range-corrected Number of Molecular I2A Photons" ;
		Nm_i2a:description = "Inverted Molecular I2A times range^2 (in m) divided by 10^6" ; 
		Nm_i2a:units = " " ;
		Nm_i2a:dpl_py_binding = "rs_inv.Nm_i2a" ;
	float Ncp(time, altitude) ;
		Ncp:long_name = "Range-corrected Number of Cross Polarized Photons" ;
		Ncp:description = "Inverted Cross Polarized times range^2 (in m) divided by 10^6" ;
		Ncp:units = " " ;
		Ncp:dpl_py_binding = "rs_inv.Ncp" ;
	float profile_Na(profile_time,altitude) ;
		profile_Na:long_name = "Range-corrected Number of Aerosol Photons" ;
		profile_Na:description = "Inverted Aerosol times range^2 (in m) divided by 10^6" ;
		profile_Na:units = " " ;
		profile_Na:dpl_py_binding = "profiles.inv.Na" ;
	float profile_Nm(profile_time,altitude) ;
		profile_Nm:long_name = "Range-corrected Number of Molecular Photons" ;
		profile_Nm:description = "Inverted Molecular times range^2 (in m) divided by 10^6" ;
		profile_Nm:units = " " ;
		profile_Nm:dpl_py_binding = "profiles.inv.Nm" ;
	float profile_Nm_i2a(profile_time,altitude) ;
		profile_Nm_i2a:long_name = "Range-corrected Number of Molecular I2A Photons" ;
		profile_Nm_i2a:description = "Inverted Molecular I2A times range^2 (in m) divided by 10^6" ;
		profile_Nm_i2a:units = " " ;
		profile_Nm_i2a:dpl_py_binding = "profiles.inv.Nm_i2a" ;
	float profile_Ncp(profile_time,altitude) ;
		profile_Ncp:long_name = "Range-corrected Number of Cross Polarized Photons" ;
		profile_Ncp:description = "Inverted Cross Polarized times range^2 (in m) divided by 10^6" ;
		profile_Ncp:units = " " ;
		profile_Ncp:dpl_py_binding = "profiles.inv.Ncp" ;
	int qc_mask(time, altitude) ;
		qc_mask:long_name = "Quality Mask" ;
		qc_mask:description = "Quality mask bitfield.  Unused bits are always high" ;
		qc_mask:missing_value = 0 ;
		qc_mask:_Unsigned = "true" ;
		qc_mask:bit_0 = "complete_mask" ;
		qc_mask:bit_0_description = "data is good.  and of bits 1-9" ;
		qc_mask:bit_1 = "lidar_ok_mask" ;
		qc_mask:bit_1_description = "lidar data is present" ;
		qc_mask:bit_2 = "lock_quality_mask" ;
		qc_mask:bit_2_description = "laser is locked to iodine filter wavelength" ;
		qc_mask:bit_3 = "seed_quality_mask" ;
		qc_mask:bit_3_description = "laser wavelength is locked to seed laser" ;
		qc_mask:bit_4 = "mol_count_snr_mask" ;
		qc_mask:bit_4_description = "molecular signal/photon counting error in molecular signal is above specified threshhold" ;
		qc_mask:bit_5 = "backscat_snr_mask" ;
		qc_mask:bit_5_description = "backscatter cross-section/photon counting error in backscatter cross-section is above specified threshhold" ;
		qc_mask:bit_6 = "mol_lost_mask" ;
		qc_mask:bit_6_description = "number of molecular photon counts is above specified threshhold" ;
		qc_mask:bit_7 = "min_backscat_mask" ;
		qc_mask:bit_7_description = "lidar backscatter cross-section is above specified threshhold" ;
		qc_mask:bit_8 = "radar_backscat_mask" ;
		qc_mask:bit_8_description = "radar backscatter cross-section is above specified threshhold" ;
		qc_mask:bit_9 = "radar_ok_mask" ;
		qc_mask:bit_9_description = "radar data is present" ;
		qc_mask:bit_10 = "aeri_ok_mask" ;
		qc_mask:bit_10_description = "aeri data is present" ;
		qc_mask:bit_11 = "aeri_qc_mask" ;
		qc_mask:bit_11_description = "aeri data has passed a quality check" ;
		qc_mask:dpl_py_binding = "rs_inv.qc_mask" ;
	float std_beta_a_backscat(time, altitude) ;
		std_beta_a_backscat:long_name = "Std dev of backscat cross section (photon counting)" ;
		std_beta_a_backscat:units = "1/(m sr)" ;
		std_beta_a_backscat:missing_value = NaNf ;
		std_beta_a_backscat:plot_scale = "logarithmic" ;
		std_beta_a_backscat:dpl_py_binding = "rs_inv.std_beta_a_backscat" ;
	short hsrl_qa_BS(time, altitude) ;
		hsrl_qa_BS:long_name = "Quality Assurance Backscatter" ;
		hsrl_qa_BS:value_NC = 0 ;
		hsrl_qa_BS:value_Good = 1 ;
		hsrl_qa_BS:value_Bad = 2 ;
		hsrl_qa_BS:value_Caution = 3 ;
		hsrl_qa_BS:dpl_py_binding = "rs_inv.qa_flags.qa_BS" ;
	short hsrl_qa_dep(time, altitude) ;
		hsrl_qa_dep:long_name = "Quality Assurance Depolarization" ;
		hsrl_qa_dep:value_NC = 0 ;
		hsrl_qa_dep:value_Good = 1 ;
		hsrl_qa_dep:value_Bad = 2 ;
		hsrl_qa_dep:value_Caution = 3 ;
		hsrl_qa_dep:dpl_py_binding = "rs_inv.qa_flags.qa_dep" ;
	short hsrl_qa_Ext(time, altitude) ;
		hsrl_qa_Ext:long_name = "Quality Assurance Extinction" ;
		hsrl_qa_Ext:value_NC = 0 ;
		hsrl_qa_Ext:value_Good = 1 ;
		hsrl_qa_Ext:value_Bad = 2 ;
		hsrl_qa_Ext:value_Caution = 3 ;
		hsrl_qa_Ext:dpl_py_binding = "rs_inv.qa_flags.qa_Ext" ;
	float rlprof_asr(time, altitude) ;
		rlprof_asr:long_name = "Raman Aerosol Scattering Ratio" ;
		rlprof_asr:units = "unitless" ;
		rlprof_asr:dpl_py_binding = "rlprofaerosol.aerosol_backscatter_ratio" ;
	float rlprof_beta(time, altitude) ;
		rlprof_beta:long_name = "Raman Beta" ;
		rlprof_beta:units = "1/(m sr)" ;
		rlprof_beta:dpl_py_binding = "rlprofaerosol.beta" ;
	float rlprof_ext_n2(time, altitude) ;
		rlprof_ext_n2:long_name = "Raman Aerosol N2 Extinction" ;
		rlprof_ext_n2:units = "1/m" ;
		rlprof_ext_n2:dpl_py_binding = "rlprofaerosol.extinction_n2" ;
	float rlprof_bscat(time, altitude) ;
		rlprof_bscat:long_name = "Raman Aerosol Backscatter Extinction" ;
		rlprof_bscat:units = "1/m" ;
		rlprof_bscat:dpl_py_binding = "rlprofaerosol.extinction_bscat" ;
	float rlprof_sa(time, altitude) ;
		rlprof_sa:long_name = "Raman Extinction to Backscatter Ratio" ;
		rlprof_sa:units = "sr" ;
		rlprof_sa:dpl_py_binding = "rlprofaerosol.extinction_to_backscatter_ratio" ;
	float rlprof_dep(time, altitude) ;
		rlprof_dep:long_name = "Raman Linear Depolarization" ;
		rlprof_dep:units = "percent" ;
		rlprof_dep:dpl_py_binding = "rlprofaerosol.linear_depol" ;

// global attributes:
        :dpl_py_template = "hsrl3_arm.cdl" ;
        :dpl_py_template_version = 20161111 ;
		:time_zone = "UTC" ;
                :code_version = "" ;
                :load_calibration_version = "" ;
                :get_internal_cal_vals_version = "" ;
                :calvals = "" ;
                :find_new_cal_times_version = "" ;
                :radiosonde_profile_version = "" ;
                :fetch_cal_version = "" ;
                :quick_cal_version = "" ;
                :processed_netcdf_version = "" ;
                :process_data_version = "" ;
                :timefill_sum_version = "" ;
                :timefill_average_version = "" ;
                :file_version = -1 ;
                :time_axis_average_mode = "obsolete" ;
                :time_axis_average_parameter = -1. ;
                :range_axis_average_parameter = -1. ;
                :featureset = -1 ;
                :featureset_version = "" ;
                :processing_parameters__qc_params__min_radar_alt = -1. ;
                :processing_parameters__qc_params__min_lidar_alt = -1. ;
                :processing_parameters__qc_params__lock_level = -1 ;
                :processing_parameters__qc_params__min_radar_dBz = -1. ;
                :processing_parameters__qc_params__backscat_snr = -1. ;
                :processing_parameters__qc_params__mol_lost = -1. ;
                :processing_parameters__qc_params__min_radar_backscat = -1. ;
                :processing_parameters__particlesettings__g_water = -1. ;
                :processing_parameters__particlesettings__h20_depol_threshold = -1. ;
                :processing_parameters__particlesettings__sigma_v = -1. ;
                :processing_parameters__particlesettings__type = "obsolete" ;
                :processing_parameters__particlesettings__alpha_ice = -1. ;
                :processing_parameters__particlesettings__p180_ice = -1. ;
                :processing_parameters__particlesettings__delta_v1 = -1. ;
                :processing_parameters__particlesettings__Dr = -1. ;
                :processing_parameters__particlesettings__g_ice = -1. ;
                :processing_parameters__particlesettings__delta_a1 = -1. ;
                :processing_parameters__particlesettings__alpha_water = -1. ;
                :processing_parameters__particlesettings__delta_v2 = -1. ;
                :processing_parameters__particlesettings__sigma_a = -1. ;
                :processing_parameters__particlesettings__delta_a2 = -1. ;
}
