netcdf out {
dimensions:
	raw_time = UNLIMITED ;
    bin_range = 0;
	time_vector = 8 ;
variables:
	int base_time ;
		base_time:string = "2006-10-23 18:19:59 UTC" ;
		base_time:long_name = "Base seconds since Unix Epoch" ;
		base_time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		base_time:dpl_py_binding = "dne" ;
	double raw_time(raw_time) ;
		time:long_name = "Raw Time" ;
		time:units = "seconds since 2006-10-23 18:19:59 UTC" ;
		time:dpl_py_binding = "rs_raw.times" ;
        time:dpl_py_type = "python_datetime" ;
	float bin_range(bin_range) ;
		bin_range:long_name = "Distance away from the lidar" ;
		bin_range:units = "meters" ;
		bin_range:dpl_py_binding = "rs_raw.msl_altitudes" ;
	float transmitted_energy(raw_time) ;
		transmitted_energy:long_name = "Transmitted Energy" ;
		transmitted_energy:units = "Joules" ;
		transmitted_energy:missing_value = 9.96920996838687e+36 ;
		transmitted_energy:dpl_py_binding = "rs_raw.transmitted_energy" ;
	int num_seeded_shots(raw_time) ;
		num_seeded_shots:long_name = "Number of Seeded Shots" ;
		num_seeded_shots:missing_value = -1 ;
		num_seeded_shots:dpl_py_binding = "rs_raw.seeded_shots" ;
	int num_shots(raw_time) ;
		num_shots:long_name = "Number of Shots" ;
		num_shots:missing_value = -1 ;
		num_shots:dpl_py_binding = "rs_raw.shot_count" ;
	float mol_cal_pulse(raw_time) ;
		mol_cal_pulse:long_name = "Molecular calibration pulse" ;
		mol_cal_pulse:description = "Sum of photon counts in the molecular channel due to light scattered with the telescope." ;
		mol_cal_pulse:units = "counts" ;
		mol_cal_pulse:missing_value = 9.96920996838687e+36 ;
		mol_cal_pulse:dpl_py_binding = "rs_raw.molecular_cal_pulse" ;
	int molecular_counts(raw_time, bin_range) ;
		molecular_counts:long_name = "Molecular Photon Counts" ;
		molecular_counts:description = "Raw counts, per averaging interval with pileup, afterpulse, and darkcount corrections applied" ;
		molecular_counts:units = "counts" ;
		molecular_counts:missing_value = -1 ;
		molecular_counts:plot_scale = "logarithmic" ;
		molecular_counts:dpl_py_binding = "rs_raw.molecular_counts" ;
	int molecular_i2a_counts(raw_time, bin_range) ;
	        molecular_i2a_counts:long_name = "Molecular I2A Photon Counts" ;
        	molecular_i2a_counts:description = "Raw counts, per averaging interval with pileup, afterpulse, and darkcount corrections applied" ;
        	molecular_i2a_counts:units = "counts" ;
         	molecular_i2a_counts:missing_value = -1 ;
        	molecular_i2a_counts:plot_scale = "logarithmic" ;
        	molecular_i2a_counts:dpl_py_binding = "rs_raw.molecular_i2a_counts" ;
	int combined_counts_lo(raw_time, bin_range) ;
		combined_counts_lo:long_name = "Low Gain Combined Photon Counts" ;
		combined_counts_lo:description = "Raw counts, per averaging interval with pileup, afterpulse, and darkcount corrections applied" ;
		combined_counts_lo:units = "counts" ;
		combined_counts_lo:missing_value = -1 ;
		combined_counts_lo:plot_scale = "logarithmic" ;
		combined_counts_lo:dpl_py_binding = "rs_raw.combined_lo_counts" ;
	int combined_counts_hi(raw_time, bin_range) ;
		combined_counts_hi:long_name = "High Gain Combined Photon Counts" ;
		combined_counts_hi:description = "Raw counts, per averaging interval with pileup, afterpulse, and darkcount corrections applied" ;
		combined_counts_hi:units = "counts" ;
		combined_counts_hi:missing_value = -1 ;
		combined_counts_hi:plot_scale = "logarithmic" ;
		combined_counts_hi:dpl_py_binding = "rs_raw.combined_hi_counts" ;
	int cross_counts(raw_time, bin_range) ;
		cross_counts:long_name = "Cross Polarized Photon Counts" ;
		cross_counts:description = "Raw counts, per averaging interval with pileup, afterpulse, and darkcount corrections applied" ;
		cross_counts:units = "counts" ;
		cross_counts:missing_value = -1 ;
		cross_counts:plot_scale = "logarithmic" ;
		cross_counts:dpl_py_binding = "rs_raw.cross_pol_counts" ;

// global attributes:
                :dpl_py_template = "segment_hsrl_raw.cdl" ;
                :dpl_py_template_version = 20140216 ;
		:time_zone = "UTC" ;
}
